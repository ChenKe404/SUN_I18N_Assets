CKT             G     2nd National Bank   第二国民银行   Abandoned Factory   废弃的工厂   Abandoned Warehouse   废弃的仓库   Abandoned Wharehouse   废弃的仓库   Adam's House   亚当的房子   Adult Visceroid   成年器官兽   Advanced Power Plant   先进发电厂   Alex-gators petshop just ahead!   前面就是鳄鱼宠物商店!   Alkaline's Battery Superstore   碱性电池超市   AlphaLightPost   灯柱   Ambrose Lounge   安布罗斯俱乐部   Ammo Crates	   弹药箱   Amphibious APC   两栖运兵车   Archer Asylum   阿切尔收容所	   Artillery	   榴弹炮   Attack Buggy	   冲锋车   Attack Cycle   突击摩托
   Automobile   汽车   Baby Visceroid   器官兽幼崽   Banshee   女妖   Barracks   兵营   Billy Bob's Harvester school   比利鲍勃的收割者学校   Blue Light Post   蓝色灯柱   Blue Tiberium Tree   蓝色泰矿树   Bostic Tower   博斯蒂克塔楼   Boxes   盒子   Bridge 1   桥梁 1   Bridge 2   桥梁 2   Bridge repair hut   修桥小屋   Business Offices   业务办公室   CABAL Obelisk   CABAL 方尖碑
   Cabal Core   CABAL 核心   Captured Commander   被俘的指挥官	   Cargo Car   货车   Carryall   吊运直升机   Chameleon Spy   变色龙间谍   Chem Lab   化学实验室   Chem Spray Infantry   毒素步兵   Chemical Missile   毒素导弹   Chemical Tank   毒素储存罐   Church   教堂	   City Hall	   市政厅   Civilian   平民   Civilian Armory   平民军械库   Civilian Array   平民设备   Civilian Hospital   平民医院   Clear Rock #1   干净的石头 #1   Clear Rock #2   干净的石头 #2   Clear Rock #3   干净的石头 #3   Clear Rock #4   干净的石头 #4   Clear Rock #5   干净的石头 #5   Component Tower   炮塔基座   Concrete Wall	   水泥墙   Connelly Court Apts.   康纳利法院酒店   Construction Yard	   建造厂   Core Defender   核心守卫   Crash 1   事故现场 1   Crash 2   事故现场 2   Crash 3   事故现场 3   Crash 4   事故现场 4   Crash 5   事故现场 5   Crate	   板条箱   Cyborg	   生化人   Cyborg Commando   生化尖兵   Cyborg Reaper   生化人收割者   D's Dog House
   D的狗屋   Daily Sun Times   每日太阳时报   Dam   水坝   Deluxe Accomodations   豪华住宿   Denzil's Last Chance Motel&   "登齐尔的最后机会"汽车旅馆   Deployed Artillery   已部署的榴弹炮   Deployed ICBM   已部署的洲际弹道导弹   Deployed Juggernaut   已部署的神像   Deployed Sensor Array   已部署的探测器   Deployed Tick Tank   已部署的蜱虫坦克   Devil's Tongue   恶魔火舌   Disc Thrower   飞盘掷弹兵	   Disruptor   声波坦克   Disruptor Turret   声波坦克炮塔   Drink YEO-CA Cola!   喝YEO-CA可乐!   Drop Pod   空投   Drop Pod Node   空投请求   Dropship	   运输船   Drum    
   E.M. Pulse   电磁脉冲
   EMP Cannon   电磁脉冲炮   Eat at Rade's Roadhouse   在雷德的路边餐厅吃饭   Elite Cadre   Elite框架   Energy Transformer	   变压器   Engineer	   工程师   Ferbie's 4 Sale   冯比斯的小卖部   Field Generator   场发生器   Fill'er Up-Pump'N'Go       Fire Storm Generator   火焰风暴
产生器   Firestorm Defense   火焰风暴
防御系统   Firestorm Wall Section   火焰风暴围墙   Fist of Nod
   NOD 之拳
   Flame Tank   火焰坦克   Flying Gas Tank   飞行油箱   Flying Tire   飞行的轮胎   Fona       GDI Hunter-Seeker   猎人导引头
   GDI Kodiak   科迪亚克   GDI Power Plant	   发电厂   GDI Tech Center   科技中心   GDI Upgrade Center   升级中心   GDI War Factory   战争工厂   Gas Pump   气泵	   Gas Pumps   气泵   Gas Station	   加油站   Gas Station Sign   加油站标志   Gate   大门   Ghost Stalker   幽灵行者   Goodie Crate   物资板条箱   Green Building   绿色建筑   Green Light Post   绿色灯柱
   Greenhouse   温室   Hamburgers $.99   汉堡 $.99   Hand Of Nod
   NOD 之手   Harpy   鸟身女妖	   Harvester	   收割者   Helipad	   停机坪   Hewitt Hair Salon   休伊特美发沙龙   Highrise Hotel   高层酒店
   Hover MLRS   悬浮火箭车   Huey the Infected Cyborg   被感染的生化人休伊   Hunter Seeker   猎人导引头   Hunting Lodge   狩猎小屋   Ice Floe   冰川   Invisible Blue Light Post   隐形蓝灯柱   Invisible Green Light Post   隐形绿灯柱   Invisible Light Post   隐形灯柱   Invisible Orange Light Post   隐形橙色灯柱   Invisible Purple Light Post   隐形紫色灯柱   Invisible Red Light Post   隐形红灯柱   Invisible Yellow Light Post   隐形黄色灯柱
   Ion Cannon	   离子炮   Ion Cannon Uplink   离子炮上行   JP       Jake McNeil   杰克·麦克尼尔   Join GDI: We save lives.   加入GDI: 我们拯救生命.
   Juggernaut   神像   Jumpjet Infantry   喷气飞行兵   Kaspm's Tiberium Warhouse   卡斯姆的泰矿仓库   Kettler's Place   凯特勒的位置   Kodiak Crash   科迪亚克坠机现场   Large Tiberium   大的泰伯利亚   Laser	   激光塔   Laser Fence Post   激光护栏   Laser Fence Section   激光围栏组   Leary Traveller Inn   利瑞旅行者旅馆   Light Infantry	   轻步兵
   Light Post   灯柱   Light Tower   灯塔   Lightner's Luxury Suites   莱特纳豪华套房   Limpet Drone   哨兵无人机   Limpet Mine   哨兵地雷   Local Inn & Lodging   当地旅馆&住宿   Local Store   当地商店
   Locomotive	   火车头   Long's Home	   隆的家
   Low Bridge   矮桥   Low Bridge End 1   矮桥桥端 1   Low Bridge End 2   矮桥桥端 2   Low Bridge End 3   矮桥桥端 3   Low Bridge End 4   矮桥桥端 4   Mammoth Mk.II   猛犸机甲   Mammoth Tank   猛犸坦克   Mammoth Tank Turret   猛犸坦克炮塔   Medic   医生   Meteorite01   陨石01   Meteorite02   陨石02   Miele Manor   米勒的庄园   Missile Launcher   导弹发射器   Missile Silo   导弹发射井   Mobile Construction Vehicle   移动工程车   Mobile EM-Pulse   移动电磁脉冲   Mobile EM-Pulse (Charged)   移动电磁脉冲(已充能)   Mobile Repair Vehicle   移动维修车   Mobile Sensor Array   移动探测器   Mobile Stealth Generator   移动隐形产生器   Mobile War Factory   移动重工   Multi-Missile   分体式导弹   Mutant	   变种人   Mutant Gun Turret   变种人碉堡   Mutant Headquarters   突变人总部   Mutant Hijacker   变种人强盗   Mutant Sergeant   变种人中士   Mutant Soldier   变种人战士   NOD Montauk	   蒙托克   NOD Power Plant	   发电厂   NOD Pyramid   NOD 金字塔	   NOD Radar   雷达   NOD Tech Center   技术中心   Negative Light Post	   负光柱   Negative Red Light	   负红光   No escape from Archer's Asylum!   无法逃离阿彻的疯人院!   Nod Hunter-Seeker   猎人导引头   Nod Spy   线人   Nod Wall   围墙   Nod War Factory   战争工厂
   North Labs   北实验室   Obelisk of Darkness   黑暗方尖碑   Obelisk of Light   光明方尖碑   Observation Tower	   观测塔   Office Building	   办公楼   Old Advanced Power Plant   老式发电厂   Old Construction Yard   老式建造厂   Old Refinery   老式采矿厂	   Old Silos   老式储存仓
   Old Temple   老式神殿   Old Weapons Factory   老式武器工厂   Only 11 miles to Zydeko's cafe!$   只有11英里到Zydeko的咖啡馆!   Orange Light Post   橙色灯柱   Orca Bomber   奥卡轰炸机   Orca Fighter   奥卡战斗机   Orca Transport   奥卡运输机   Oxanna   奥克斯安娜   Palette	   调色板   Pannullo Hacienda   潘努洛财政部   Pannullo's hacienda es bueno   潘努洛的财政状况很好   Panullo Hacienda   潘努洛的庄园   Passenger Car   乘客车厢   Pavement   强化地面   Pickup Truck   皮卡   Port-A-Shack	   小板房   Port-A-Shack Deluxe   豪华的小板房   Power Turbine   动力涡轮机   Purple Light Post   紫色灯柱   Pyramid	   金字塔   RPG Upgrade   榴弹   Radar   雷达   Radar Relay	   雷达站   Rade's Roadhouse   雷德的路边酒店   Railroad Bridge 1
   铁路桥1   Railroad Bridge 2
   铁路桥2   Recreational Vehicle	   休闲车   Red Light Post   红色灯柱   Regulator Station	   调节站   Relay Station	   中继站   Research Facility   研究设施   Rocket Infantry	   火箭兵   Rooms $29 a nite   房间 $29 每晚   SAM Upgrade   防空导弹   Sam   萨姆飞弹   Sand Rock #1
   1号砂岩   Sand Rock #2
   2号砂岩   Sand Rock #3
   3号砂岩   Sand Rock #4
   4号砂岩   Sand Rock #5
   5号砂岩   Sandbags   沙袋   Sandberg and Son's   桑德伯格父子公司
   School Bus   校车   Scrap Metal Debris   废金属碎片
   Scrin Ship   思金飞船   Seeker Control   猎人导引头   Service Depot	   维修坪   Slavick   斯拉维克   Solar Panel   太阳能电池板
   South Labs   南实验室   Stealth Generator   隐形产生器   Stealth Tank   隐形坦克   Stop in at Hewitt's hair salon'   在休伊特的美发沙龙稍作停留   Subterranean APC   钻地运兵车   Subterranean Dwelling   地下住宅   T.V. Station	   电视塔   TacticX games rock!   战术X游戏摇滚!   Tall's Residence   塔尔的住宅
   Technician	   技术员   Temp Housing   临时住房   Temple of NOD   神殿   The Projects   项目   Threat Rating Node   威胁等级节点   Tiberian Fiend   泰伯野兽   Tiberian Sun - Firestorm!   泰伯利亚之日 - 火焰风暴,   Tiberian Sun -- Official Rules of Engagement(   泰伯利亚之日 -- 官方交战规则   Tiberium   泰伯利亚   Tiberium (Blue)   泰伯利亚 (蓝色)   Tiberium (Green)   泰伯利亚 (绿色)   Tiberium (Large)   泰伯利亚 (大)   Tiberium Aboreus       Tiberium Cruentus   泰伯利亚 Cruentus   Tiberium Floater   泰伯利亚漂浮物   Tiberium Refinery   泰矿精炼厂   Tiberium Riparius       Tiberium Silo   泰矿储存仓   Tiberium Tree   泰伯利亚树   Tiberium Veins   泰伯利亚脉络   Tiberium Vinifera   泰伯利亚葡萄   Tiberium Waste Facility   泰矿物质回收厂   TiberiumCrystal01   泰伯利亚水晶01   TiberiumCrystal02   泰伯利亚水晶02   TiberiumShard   泰伯利亚碎片	   Tick Tank   蜱虫坦克   Titan   泰坦   Toxin Soldier   毒素步兵   Track EW	   轨道 EW   Track NS	   轨道 NS
   Track NeSw   轨道 NeSw
   Track NwSe   轨道 NwSe	   Train Car   火车车厢   Train Station	   火车站   Train Tracks   火车轨道   Tratos   特拉托斯   Tree   树   Truck   卡车   Truck (loaded)   卡车(装载)   Umagon	   乌玛贡   Urban Housing   城市住房   Urban Storefront   城市店面   Vega's Pyramid   维加的金字塔   Veinhole Monster   脉络孔怪物   Veinhole Monster Dummy   脉络孔假人   Veinhole Tree   脉络孔树   Visit Scenic Las Vegas   游览拉斯维加斯风景区   Vulcan Cannon   火神机枪   WS Logging Company   WS测井公司   WW Surf and Turf hits the spot!   WW Surf and Turf精彩纷呈!   Water Purifier   污水处理厂
   Water Tank   水箱
   Waystation	   中转站
   Weed Eater	   回收者   Westwood Stock Exchange   Westwood证券交易所	   Wolverine   狼獾   YEO-CA Cola Corp.   YEO-CA 可乐公司   Yee's Discount Liquor   易的折扣酒吧   Yellow Light Post   黄色灯柱battle       (   Act 1: GDI Campaign - Desperate Measures   GDI战役 - 亡命之计3   Act 2: Brotherhood of Nod Campaign - From the Ashes!   Nod兄弟会战役 - 灰烬重生*   Brotherhood of Nod Campaign - Deus ex Kane'   Nod兄弟会战役 - 凯恩杀出重围$   GDI Campaign - Evolutionary Response   GDI战役 - 进化反应
fs_mission    $   �  CABAL has betrayed us all. GDI and perhaps the Earth itself are doomed unless we can fall back and regroup in time to send for help. The first priority is to deliver Dr. Boudreau to the nearby GDI outpost for immediate evacuation. Once safe, she will call for additional reinforcements.@END TRANSMISSION.@@First Objective: Escort Dr. Boudreau to the GDI outpost for immediate evacuation.@@Second Objective: Fortify this outpost and destroy CABAL’s base.�  CABAL背叛了我们所有人. GDI, 甚至整个地球都要完蛋了, 不过只要我们能够及时撤退就还有机会东山再起. 首要任务是将 Boudreau 博士护送至附近的GDI前哨站进行紧急撤离. 一旦她安全, 她将呼叫增援部队. @通讯结束.@@目标一: 护送 Boudreau 博士前往GDI前哨站以便紧急撤离. @@目标二: 加固前哨站并摧毁CABAL的基地.#  CABAL has betrayed us all. We must escape and regroup in order to repay him for his treachery. There is an abandoned airfield nearby; if we can reach it, we have a chance. Once there, we must repair the array to contact our forces and call for an immediate evacuation. We have no information or tactical support now that CABAL has gone rogue.@DATA LINK CLOSED.@@First Objective: Evade CABAL's forces and find the abandoned airfield.@@Second Objective: Repair the array to call for an immediate evacuation.@@Third Objective: Retreat to the Montauk.�  CABAL背叛了我们所有人. 我们必须撤离并重整队伍, 回头再清算他的背叛行为. 附近有一座废弃的机场, 如果我们能抵达那里, 就还有一线生机. 到达后, 我们必须修复通讯设备以向我方部队发送撤离请求. 如今CABAL已叛变, 我们没有任何情报或战术上的支援. @数据链接关闭.@@目标一: 避开CABAL的部队并找到废弃机场. @@目标二: 修复通讯设备以请求撤离. @@目标三: 撤退到蒙托克.�  CABAL's core has been disassembled and is in the hands of GDI. With the Brotherhood in a state of disarray it is essential to get CABAL back online. Locate and retrieve the three pieces of the core without alerting the local GDI forces. Remaining silent is the only hope for a successful operation.@DATA LINK CLOSED.@@First Objective: Infiltrate the GDI base.@@Second Objective: Locate the three pieces of CABAL's core.@@@Third Objective: Return to the drop zone for immediate retrieval and evacuation.}  CABAL的核心已被拆解, 目前掌握在GDI手中. 随着兄弟会陷入混乱状态, 恢复CABAL的运行至关重要. 在不惊动当地GDI部队的情况下定位并取回三块核心组件. 保持隐蔽是行动成功的唯一手段. @数据链接关闭.@@目标一: 潜入GDI基地。@@目标二: 找到CABAL核心的三块组件. @@@目标三: 返回空投区域并撤离.J  CABAL’s core is believed to be in this area. Using an engineer, infiltrate and capture the core. Cut off enemy reinforcements by destroying the two bridges that supply this base. Nod is utilizing self-powered laser fencing to protect the core from intruders. Disable this fencing by capturing the appropriate command stations using local civilian technicians. Once inside, neutralize any remaining defense systems guarding the core.@END TRANSMISSION.@@First Objective: Destroy the two bridges to stem the flow of reinforcements.@@Second Objective: Infiltrate and capture CABAL's core.�  据情报, CABAL的核心位于该区域. 利用工程师渗透并夺取该核心. 通过摧毁连接该基地的两座桥梁来切断敌方增援. Nod正在使用自供能的激光围栏来防止入侵者接近核心. 通过让当地平民技术员占领相关指挥站来关闭这些围栏. 一旦进入, 清除核心周围所有的防御系统. @通讯结束.@@目标一: 摧毁两座桥梁以阻止敌方增援. @@目标二: 渗透并夺取CABAL的核心.   GDI 01:Recover the Tacitus   GDI 01: 取回塔西佗   GDI 02:Party Crashers   GDI 02: 派对破坏者   GDI 03:Quell the Civilian Riot   GDI 03: 镇压平民暴动   GDI 04: In the Box   GDI 04: 在盒子里   GDI 05: Dogma Day Afternoon   GDI 05: 礼拜日的下午   GDI 06:Escape from CABAL   GDI 06: 从CABAL撤离   GDI 07: The Cyborgs are Coming   GDI 07: 生化人来了   GDI 08:Factory Recall   GDI 08: 工厂召回   GDI 09:Core of the Problem   GDI 09: 问题的核心B  GDI scientists have reprogrammed a NOD cyborg and have implanted a virus designed for release into CABAL's communications network. The cyborg must be inserted into CABAL's defensive outpost for the virus to take effect. CABAL is aware of this operation and will do anything to prevent it. Establish your base quickly before CABAL can fortify his position.@END TRANSMISSION.@@First Objective: Insert the infected cyborg into the defensive outpost's network center.@@Second Objective: Destroy the cyborg manufacturing facility.@Third Objective: Destroy all remaining CABAL forces.�  GDI科学家重写了一个Nod生化人的程序, 并植入了一种用于释放到CABAL通讯网络中的病毒. 你必须将这个生化人送入CABAL的防御前哨站, 病毒才能生效. CABAL已经得知这次行动, 会不择手段地阻止你. 在CABAL加固防御之前, 迅速建立你的基地. @通讯结束.@@目标一: 将感染病毒的生化人送入前哨站的网络中心. @@目标二: 摧毁生化人制造设施. @目标三: 消灭所有剩余的CABAL部队.   NOD 01:Operation Reboot   NOD 01: 操作重新启动   NOD 02:Seeds of Destruction   NOD 02: 毁灭的种子   NOD 03:Tratos’ Final Act   NOD 03: 特拉托斯的终幕   NOD 04:Mutant Extermination   NOD 04: 变种人灭绝   NOD 05:Escape from CABAL   NOD 05: 逃离CABAL   NOD 06: The Needs of the Many!   NOD 06: 许多人的需求!   NOD 07: Determined Retribution   NOD 07: 坚决的惩罚   NOD 08: Harvester Hunting   NOD 08: 收割者猎人   NOD 09:Core of the Problem   NOD 09: 问题的核心7  Prior to our main assault on CABAL, we need to slow down his production capabilities. CABAL is harvesting Tiberium heavily in Eastern Africa. Proceed there and eliminate CABAL's harvesting facilities. Our forces are scattered at this time and we can only afford to provide you with a small strike force.@@Use the new Fist of Nod mobile production facility to build up an effective strike force and crush them.@DATA LINK CLOSED.@@First Objective: Save the Civilians and their town from CABAL's siege.@@Second Objective: Disrupt and prevent CABAL's Tiberium harvesting.�  在我们对CABAL发动主攻之前, 必须先削弱他的生产能力. CABAL正在非洲东部大规模开采泰伯利亚. 前往该地区并摧毁CABAL的采集设施. 目前我方兵力分散, 只能为你提供一支小型突击部队. @@使用新的Nod之拳移动工厂来组建有效的打击力量并将其摧毁. @数据链接关闭.@@目标一: 从CABAL的围攻中解救平民及其城镇. @@目标二: 破坏并阻止CABAL采集泰伯利亚.

�  Scorched earth, plain and simple. Locate and destroy all cybernetic forces in the area. The base has a web of laser fences protecting it and CABAL's computer core.@DATA LINK CLOSED.@@First Objective: Repair the bridges to allow for reinforcements.@@Second Objective: Capture the command station to shut down the laser fencing surrounding CABAL's core.@@Third Objective: Destroy CABAL's base and all defenses.F  焦土战略, 找到并消灭该区域内的所有生化人部队. 该基地布满了激光围栏, 用以保护CABAL的计算核心.@数据链接关闭.@@目标一: 修复桥梁以便增援部队通行. @@目标二: 占领指挥站以关闭围绕CABAL核心的激光围栏. @@目标三: 摧毁CABAL的基地及其所有防御.�  Since CABAL has turned on us we are suffering a communications blackout. We are forced to try and obtain GDI's EVA technology. There is a small GDI airbase in this sector. Get your engineer into their radar facility to steal an EVA unit. Create a distraction to occupy GDI air units while you steal the EVA unit.@@We also have a new unit for you: the Mobile Stealth Generator is now operational. Use it wisely.@DATA LINK CLOSED.@@First Objective: Reconnoiter the area to find the GDI base and civilian towns.@@Second Objective: Create distractions to draw away the GDI base's air support.@@Third Objective: Get an engineer into GDI's radar facility to steal the EVA unit.�  由于CABAL的背叛, 我们的通讯中断了. 我们被迫试图获取GDI的EVA技术. 这个区域有一个小型GDI空军基地, 派遣你的工程师潜入雷达设施, 制造干扰以牵制GDI空中单位, 同时窃取EVA单元. @@我们为你准备了一种新单位: 移动隐形发生器. @数据链接关闭.@@目标一: 侦察区域, 找到GDI基地及平民城镇. @@目标二: 制造干扰, 牵制GDI基地的空中支援.@@目标三: 派工程师潜入GDI雷达设施, 窃取EVA单元.~  The Kodiak was lost en route to the Philadelphia. We believe it has crashed somewhere in the area. The Kodiak was carrying the recently recovered Tacitus when it went down. Take a small team and locate the crash site and determine if the Kodiak can be repaired. Recover the Tacitus at all costs. Be advised, there are reports that NOD forces and hostile Tiberian life forms have been sighted in the area. The ion storm is still in full force, so advanced units cannot be used.@END TRANSMISSION.@@First Objective: Find the Kodiak and determine if it can be salvaged.@@Second Objective: Recover the Tacitus and return it to the pickup zone.  科迪亚克号在前往费城的途中失联. 我们知道它在该区域某处坠毁了. 科迪亚克号坠毁时携带了最近回收的塔西佗. 带领一支小队找到坠毁地点, 评估科迪亚克是否还能修复. 无论代价如何, 都要回收塔西佗. 注意, 有报告称该区域出现了Nod部队和敌对的泰伯生命体. 离子风暴仍在持续发生, 故无法使用高级单位. @通讯结束.@@目标一: 找到科迪亚克并评估是否可回收. @@目标二: 回收塔西佗并送回接收区.�  The death of Tratos has caused open revolt among the mutant population. They believe the local food and water supplies have been poisoned and are attacking the local supply depot. This has aggravated civilian tensions in the area causing armed conflict between the two factions.@@Deploy your squad and quell the rioting.  Prevent casualties and damage on BOTH sides of the conflict. To this end we have equipped your infantry with non-lethal weaponry. In addition, you must prevent the destruction of the depot as it supplies all of the relocated civilians and mutants in the area.@END TRANSMISSION.@@First Objective: Neutralize the four riot leaders without killing any of the civilians or mutants.@@Second Objective: Prevent the Supply Depot from being destroyed.X  特拉托斯的死引发了变种人群体的公开暴动. 他们认为当地的食物和水源被下了毒, 正在攻击当地的补给仓库. 这加剧了该地区民众的紧张局势, 导致双方发生武装冲突. @@派遣你的队伍平息骚乱. 防止冲突双方人员伤亡和财产损失. 为此, 我们为你的步兵配备了非致命武器. 此外, 你必须防止补给仓库被毁, 因为它为该地区所有被安置的平民和变种人提供补给.@通讯结束.@@目标一: 制服四名暴乱头目, 且不得伤害任何平民或变种人.@@目标二: 防止补给仓库被毁.  The first step in our Tiberium evolution requires the fertilization of the land with new indigenous life forms. We will use this new life to educate those who wish to interfere with its progress. Locate and repair the bridge leading to the Genesis Pit before using the Toxin Soldiers to "persuade" the nearby civilians to aid us in our cause.@DATA LINK CLOSED.@@First Objective: Remain hidden from the GDI forces in the area.@@Second Objective: Use drugged civilians to lure life forms out of the Genesis Pit to cleanse the region.�  泰伯利亚进化的第一步是用新的本土生命体来肥沃土地. 我们将利用这些新的生命体"教育"那些试图干涉其进展的人. 在使用毒素步兵"说服"附近平民协助我们之前, 先找到并修复通往创世纪坑的桥梁. @数据链接关闭.@@目标一: 避免被GDI部队发现.@@目标二: 利用被下药的平民诱导生命体走出创世纪坑, 以净化该区域.<  The mutant vermin have once again made themselves known to us. They have stolen the Tacitus that I...we have worked so hard to obtain. If Kane's vision is to be fulfilled, we must find the mutant encampment and recover the Tacitus. Once it is safely removed, terminate any mutants who decide to remain in the area. Perhaps this will teach them not to interfere with us ever again.@DATA LINK CLOSED.@@First Objective: Locate the mutant encampment.@@Second Objective: Recover the Tacitus and return it to the drop zone.@@Third Objective: Destroy all remaining mutant forces.�  变种害兽再次现身. 他们偷走了我...我们费尽心力获得的塔西佗. 若要实现凯恩的愿景, 我们必须找到变种人营地并夺回塔西佗. 安全取回塔西佗后, 消灭任何选择留在该区域的变种人. 也许这能教训他们以后不要再来挑衅我们. @数据链接关闭.@@目标一: 找到变种人营地. @@目标二: 夺回塔西佗并送回空投区. @@目标三: 消灭所有剩余的变种人部队.9  The second piece of the Tacitus is rumored to be held inside an ancient temple outside of La Paz, Bolivia. Ghoststalker and one of our archaeologists will assist you in locating the temple and retrieving the Tacitus.@We also have a new unit for you to test: it's called the Juggernaut and is our new long-range artillery unit. Be advised: this area is completely uncharted.@END TRANSMISSION.@@First Objective: Reconnoiter the area and identify the Temple of the Tacitus.@@Second Objective: Recover the Tacitus from the temple and proceed to the designated airlift zone.�  据传塔西佗的第二块碎片被藏在玻利维亚拉巴斯外的一座古老神殿中. 幽灵行者和我们的考古学家将协助你找到该神殿并取回塔西佗. @我们还为你准备了一种新单位供测试: 它被称为"巨兽", 是我们的新型远程火炮单位. 请注意: 该区域是完全未知的. @通讯结束.@@目标一: 侦察区域并确认塔西佗神殿的位置.@@目标二: 从神殿中回收塔西佗并前往空投区.�  This is it Commander! Take out CABAL fast and hard: No mercy and no surrender. Find a way to get inside his defenses and take out the core. GDI forces are distracting CABAL and now is the perfect time to crush CABAL once and for all.@DATA LINK CLOSED.@@First Objective: Build your base and survive the initial onslaught from CABAL.@@Second Objective: Capture the 3 control stations to shut down the laser fences and firestorm defense system protecting CABAL.@@Third Objective: Destroy CABAL’s core.�  就是现在, 指挥官! 猛烈地痛击CABAL, 毫不留情, 绝不手软.找到进入防线的途径, 摧毁CABAL核心. GDI部队正在牵制CABAL, 现在正是彻底粉碎他的最佳时机. @数据链接关闭.@@目标一: 建立基地并挺过CABAL的首次猛攻. @@目标二: 占领3个控制站以关闭保护CABAL的激光围栏和火风暴防御系统. @@目标三: 摧毁CABAL的核心.�  We have lost communication with a small civilian settlement nearby. Incoming messages from our remote base indicate an attack from unidentified life forms. Investigate these sightings and protect the civilians at all costs. Escort as many civilians as possible to the pickup zone for immediate evacuation.@END TRANSMISSION.@@First Objective: Protect the small clusters of civilians and escort them to the designated airlift zone.@@Second Objective: Defend the base from attacks until reinforcements arrive.q  我们与附近一个小型平民定居点失去了联系. 远程基地传来消息, 称受到不明生命体的袭击. 调查这些目击事件, 并不惜一切代价保护平民. 护送尽可能多的平民到接送区进行紧急撤离.@通讯结束.@@目标一: 保护小型平民聚居点并护送他们到指定区域. @@目标二: 在援军到达前防御基地.`  We have lost communication with our base outside of Trondheim. Scout the area and determine the cause of this interruption. We have no tactical data on CABAL's forces in that area and we need information.@END TRANSMISSION.@@First Objective: Warn the local civilians of the CABAL threat.@@Second Objective: Establish a base and destroy CABAL’s forces.   我们与特隆赫姆外的基地失去了联系. 侦察该区域, 查明通讯中断的原因. 另外, 我们没有该区域内CABAL部队的情报. @通讯结束.@@目标一: 警告当地平民CABAL的威胁.@@目标二: 建立基地并摧毁CABAL部队.  We've tracked down CABAL and are ready to engage his forces on all fronts. This is an all-out assault. Nod forces have reluctantly agreed to a temporary cease-fire and are launching their own simultaneous offensive against CABAL. Destruction of the core is essential to our victory.@END TRANSMISSION.@@First Objective: Build a base and repel initial attacks.@@Second Objective: Capture the 3 control stations to shut down the laser fences and firestorm defense system protecting CABAL.@@Third Objective: Destroy CABAL’s Core.@�  我们已追踪到CABAL, 准备在各个战线发起攻击. 这是一场全面进攻. Nod部队勉强同意暂时停火, 并对CABAL发起协同进攻. 摧毁核心对我们的胜利至关重要. @通讯结束.@@目标一: 建立基地并抵御初期攻击. @@目标二: 占领3个控制站以关闭保护CABAL的激光围栏和火风暴防御系统.@@目标三: 摧毁CABAL的核心.@C  While GDI forces have been diverted to defend civilians, you are to lead an elite strike force to assassinate the mutant leader Tratos. Our new limpet mines will help you locate Tratos within his fortified base. Once located you must devise a way to reach him. GDI will have considerable protection for Tratos as he is their last hope at countering the Tiberium onslaught. Destroying their power supply should neutralize the firestorm defense system, and an effective air strike should deal with the sensor arrays.@@Do not fail: this mission is integral to the future of the Brotherhood of Nod.@DATA LINK CLOSED.@@First Objective: Attach limpet mines to GDI units to penetrate the base and locate Tratos.@@Second Objective: Deactivate the firestorm defense system and neutralize the sensor arrays.@@Third Objective: Assassinate Tratos.�  当GDI部队被调往保护平民时, 你将率领一支精英突击队刺杀变种人首领特拉托斯. 我们新型的磁吸地雷将帮助你在其设防基地内定位特拉托斯. 找到目标后, 你必须想办法接近他. GDI将为特拉托斯提供强力保护, 因为他是抵御泰伯利亚攻击的最后希望. 摧毁其电力来源应该可以使火风暴防御系统失效, 空袭则应该能摧毁传感器阵列. @@绝不能失败: 此任务关系兄弟会的未来. @数据链接关闭.@@目标一: 将磁吸地雷附着于GDI单位, 以渗透基地并定位特拉托斯.@@目标二: 关闭火风暴防御系统并摧毁传感器阵列. @@目标三: 刺杀特拉托斯.fs_tutorial    �      "Temple of Thunder"   "雷光神殿"   "Temple of Time"   "时光神殿"   "Temple of the Tacitus"   "塔西佗神殿"'   ****BATTLEFIELD CONTROL ESTABLISHED****   ****作战控制已连接****:   ****ESTABLISHING BATTLEFIELD CONTROL****..........Standby!-   ****作战控制连接中****  ... 请稍候!+   A piece of CABAL's core has been recovered.&   CABAL核心的一部分已经被找到   ARCHAEOLOGIST killed!   考古学家被杀了!   Aircraft approaching.   飞机正在接近=   Archaeologist: Command, this is Valdez, I've got the Tacitus!C   考古学家: 指挥部, 我是瓦尔迪兹, 我找到塔西佗了!3   Archaeologist: The Hieroglyphs on this temple read:6   考古学家: 神殿上的象形文字是这样写的:v   CABAAL: During the Ion Storm their Radar/Communications will be down. Now is the opportune time to hit them before thec   CABAL: 离子风暴期间, 他们的雷达/通讯将会中断. 现在正是打击他们的好时机3   CABAAL: GDI Communications have been reestablished.   CABAL: GDI通讯已经重建   CABAL on-line...   CABAL 上线...8   CABAL: Arrays have been destroyed, sensors are now down.0   CABAL: 阵列已被摧毁, 传感器也失灵了0   CABAL: SAM sites destroyed.  Air power incoming.3   CABAL: 萨姆飞弹基地已被摧毁. 空军来袭L   CABAL: The capture of 6 power plants will shut down the Firestorm Generator.;   CABAL: 占领6座发电厂就能关闭火焰风暴发生器C   CABAL: You have been detected, Tratos is escaping by air transport.?   CABAL: 你们被发现了, 特拉托斯正在乘坐飞机逃跑+   CABAL: You have failed, Tratos has escaped.-   CABAL: 你们失败了, 特拉托斯逃走了   CIVILIAN CASUALTY TOO HIGH!   平民伤亡太高!
   CIVILIANS.   平民;   Cabaal: Establish a foothold on the far side of this bridge1   CABAL: 在这座桥的另一边建立一个防线;   Cabaal: Hassan's Base has been alerted. Attack is imminent.8   CABAL: 哈桑基地已经收到警报.攻击迫在眉睫)   Cabaal: MCV has arrived to the southeast.   CABAL: MCV已经到达东南方�   Cabal: Find and capture the train station before Umagon arrives. If she manages to make it onto a train then destroy it before she can escape.x   CABAL: 在乌玛贡到达之前找到并占领火车站. 如果她成功登上了火车那就在她逃脱之前摧毁它B   Cabal: General Vega, the generators are online.  SAM sites active.J   CABAL: 维加将军, 发生器已经启动. 萨姆飞弹发射台已激活M   Cabal: General Vega, the secondary generators will come online in 20 minutes.>   CABAL: 维加将军, 第二台发生器将在20分钟内启动<   Cabal: Power plant eliminated. 1 left to capture or destroy.+   CABAL: 发电厂已被清除, 还剩余1座<   Cabal: Power plant eliminated. 2 left to capture or destroy.+   CABAL: 发电厂已被清除, 还剩余2座<   Cabal: Power plant eliminated. 3 left to capture or destroy.+   CABAL: 发电厂已被清除, 还剩余3座<   Cabal: Power plant eliminated. 4 left to capture or destroy.+   CABAL: 发电厂已被清除, 还剩余4座<   Cabal: Power plant eliminated. 5 left to capture or destroy.+   CABAL: 发电厂已被清除, 还剩余5座!   Can I offer you a tasty beverage?   要来杯可口的饮料吗?   Can anyone help us?   有人能帮帮我们吗?$   Civilian: HELP! We are under attack!&   平民: 救命! 我们受到攻击了!7   Civilian: MAYDAY! MAYDAY! We are currently under siege.*   平民: 求救! 求救! 我们被包围了/   Cult Member: Welcome Traveler! Have you come to2   邪教成员: 欢迎旅行者! 你醒过来了吗?8   Cyborg Commando online. Retaliation protocols initiated.&   生化尖兵上线. 报复协议启动k   EVA: Enemy Bridges may allow for unit reinforcement. Their destruction would be beneficial to this mission.R   EVA: 敌人的桥梁可能允许部队增援. 摧毁它们将有利于这次任务�   EVA: Locating fence technicians may help in shutting down the laser fencing. Their probable location is within a civilian outpost to the north.m   EVA: 找到围栏技术人员可能有助于关闭激光围栏. 他们可能在北边的一个平民前哨站M   EVA: Nod has aquired the Tacitus.  Recover it and return it to the drop zone.=   EVA: Nod盗取了塔西佗, 把它夺回来并带到撤离点3   EVA: Proceed to the base and secure it from attack.#   EVA: 去基地保护它不受攻击E   Escort the civilians to the ORCA transports for an immediate airlift.-   护送平民到奥卡运输机并立即撤离Z   First Objective: Attach limpet mines to GDI units to penetrate the base and locate Tratos.P   目标一: 在GDI单位上安装帽贝地雷以穿透基地并找到特拉托斯3   First Objective: Destroy all of CABAL's HARVESTERS,%   目标一: 摧毁CABAL所有的矿车=   First Objective: Find and evacuate any civilians in the area.,   目标一: 找到并疏散该地区的平民!   First Objective: Find the Kodiak.   目标一: 找到科迪亚克Y   First Objective: Get an Engineer into the Temple of Nod to retrieve part of CABAL's core.C   目标一: 让一名工程师进入Nod神殿取回部分CABAL核心I   First Objective: Get the infected Cyborg into the communications network.5   目标一: 让受感染的生化人进入通讯网络(   First Objective: Get to the GDI outpost.   目标一: 到达GDI哨所(   First Objective: Locate the Mutant base.    目标一: 找到变种人基地/   First Objective: Locate the abandoned airfield.    目标一: 找到废弃的机场@   First Objective: Neutralize (do not kill) the four riot leaders.1   目标一: 中立(不杀死)四个暴乱领导人?   First Objective: Remain hidden from the GDI forces in the area.&   目标一: 在该地区躲避GDI部队/   First Objective: Use your commander to warn the)   目标一: 使用你的指挥官警告敌4   GDI Command: Roger that Valdez, Transport is dusting<   GDI指挥部: 收到, 瓦尔迪兹号, 运输机正在前往2   GDI Command: We are providing you with a new unit,2   GDI指挥部: 我们将为你提供一支新部队4   GDI Commander: Arm Yourselves! CABAL is conscripting-   GDI指挥官: 武装起来! CABAL正在征兵*   GDI Commander: Attention Mutants! CABAL is'   GDI指挥官: 变种人注意! CABAL是*   GDI Commander: Be warned! CABAL has set up*   GDI指挥官: 小心! CABAL已经初始化1   GDI Commander: My God! CABAL is taking prisoners?1   GDI指挥官: 我的老天: CABAL正在抓人质?,   GDI Commander: People of Trondheim, you must1   GDI指挥官: 特隆赫姆的人民, 你们必须'   GDI Commander: This must be the base...&   GDI指挥官: 这肯定就是基地...   GDI Commander: What the...!?   GDI指挥官: 什么鬼!?=   GDI Soldier: Sir, these laser posts are stronger then normal.@   GDI士兵: 长官, 这些激光塔感觉比普通的还要厉害   GDI forces are near!   GDI部队就在附近!   GDI has detected your presence.   GDI侦测到你的存在"   GDI is moving a piece of the core.   GDI是一块移动的核心1   Get to the pick up zone for immediate evacuation!   到集结地立即撤离!)   Get your ENGINEER to the evacuation zone.   让你的工程师去撤离区'   Get your people to the evacuation zone.   让你的人去撤离区   HARVESTER for your troubles.    0   Here Commander, please take these two DISRUPTERS1   这里, 指挥官, 请带上这两个声波坦克   I am the power and the glory!"   我就是力量和荣耀的化身!1   Intercept the core piece before it is trasported.'   在核心部件被运走之前拦截它   Jebediah Smith?       Join us!   加入我们!?   Lead the Tiberium life forms to the GDI/civilian occupied area.+   把泰矿生命体带到GDI/平民占领区   MCV and good luck.   基地车并祝你好运&   Mayor: Yes, yes. I will see to it that'   市长: 是的, 是的. 我会注意的   Montauk Destroyed!   已摧毁蒙托克!7   Mutant Guard: Halt, and prepare for vehicle inspection!+   变种人守卫:停车, 准备车辆检查!,   Mutant Guard: It's bugged... Destroy it now!3   变种人守卫: 它被窃听了...赶快毁了它!,   Mutant Guard: Okay, looks good.  Head on in.1   变种人守卫:好的, 看起来不错.头朝里$   Mutant: Understood Blunt!  Take this#   变种人:明白直率!尝尝这个#   Mutant: We've got you now Nod scum!%   变种人:我们抓到你了, 蠢货!1   Nod General: Commander, GDI command has requested   指挥官, GDI命令已请求+   Nod General: Forget the Civilians, they are(   Nod将军: 忘掉平民吧, 他们就是/   Nod General: Well done, Commander.  GDI Command%   Nod将军:干得好, 司令.GDI命令2   Nod General: Well done, Commander.  Reinforcements(   Nod将军:干得好, 司令.增援部队(   Nod Soldier: Let's get those harvesters!$   Nod士兵: 我们去找那些矿车!(   Nod Soldier: This should be easy enough.   Nod士兵:这应该很容易3   Nod: CABAL forces are attacking! Evacuate the base!)   Nod:CABAL部队正在进攻!撤离基地!6   Now get an engineer over here to fix this bridge and I)   现在找个工程师来修这座桥, 我.   Objective Four: Destroy the research facility.   目标四: 摧毁研究设施\   Objective One: Build a Tiberium Refinery and begin harvesting the Tiberium to the southeast.I   目标一: 建造一座泰矿精炼厂, 并开始在东南方开采泰矿9   Objective One: Capture Hassan's T.V. station to the east.)   目标一: 占领东部哈桑的电视台:   Objective One: Capture the GDI base before McNeil arrives.5   目标一: 在麦克尼尔到达之前占领GDI基地h   Objective One: Capture the remaining GDI structures within this base to build a force to capture Tratos.R   目标一: 占领基地内剩余的GDI建筑, 组建一支部队占领特拉托斯K   Objective One: Contact the mutants - try searching near the local hospital.G   目标一: 与变种人取得联系 - 尝试在当地医院附近搜索:   Objective One: Deploy the ICBM launchers near the beacons.;   目标一: 在信标附近部署洲际弹道导弹发射器+   Objective One: Destroy Nod missile complex.    目标一: 摧毁Nod导弹基地3   Objective One: Destroy all of Hassan's elite guard.,   目标一: 摧毁哈桑的所有精锐卫队'   Objective One: Destroy the supply base.   目标一: 摧毁补给基地D   Objective One: Establish a base and build a Tiberium Waste Facility.&   目标一: 建造泰矿物质回收厂    Objective One: Establish a base.   目标一: 建立基地&   Objective One: Find and rescue Oxanna.)   目标一: 找到并营救奥克斯安娜@   Objective One: Infiltrate the GDI Communication Upgrade Centers.    目标一: 渗透GDI通信中心+   Objective One: Locate and free the mutants.#   目标一: 找到并释放变种人0   Objective One: Locate and secure the crash site.&   目标一: 找到并保护坠机现场:   Objective One: Locate the abandoned Nod base to the north.2   目标一: 将废弃的诺德基地定位在北部P   Objective One: Locate the crashed UFO and retrieve Kane's artifacts from inside.L   目标一: 找到坠毁的不明飞行物, 并从里面取回凯恩的文物,   Objective One: Locate the old Temple of Nod.   目标一: 寻找Nod神庙'   Objective One: Locate the toxin trucks.&   目标一: 找到运送毒素的卡车4   Objective One: Plant C4 on all ten Nod power plants..   目标一: 在所有十座Nod发电厂安装C4/   Objective One: Protect the Kodiak at all costs./   目标一: 不惜一切代价保护科迪亚克7   Objective One: Stop the launch of the Tiberium Missile.#   目标一: 阻止泰矿导弹发射4   Objective Three: Destroy all Nod forces in the area.)   目标三: 摧毁区域内所有Nod部队(   Objective Three: Destroy all Nod forces.    目标三: 摧毁所有Nod部队A   Objective Three: Get McNeil into the APC at the extraction point./   目的三: 在撤离点让麦克尼尔进入APC;   Objective Three: Locate the research facility to the north.&   目标三: 找到北方的研究设施8   Objective Two: Build a Barracks to create more infantry.7   目标二: 建立一个兵营, 以培养更多的步兵'   Objective Two: Build the Temple of Nod.   目标二: 建造Nod神殿-   Objective Two: Capture Nod Technology Center.#   目标二: 捕捉结节技术中心9   Objective Two: Clear both ends of the tunnel to the west.&   目标二: 清除隧道西面的两端0   Objective Two: Commandeer a transport to escape.#   目标二: 征用运输工具撤离1   Objective Two: Destroy Hassan's elite guard base.,   目标二: 摧毁哈桑的精英卫队基地&   Objective Two: Destroy all Nod forces.    目标二: 摧毁所有Nod部队.   Objective Two: Destroy all five Nod SAM sites.0   目标二: 摧毁所有五个防空导弹基地.$   Objective Two: Destroy the GDI base.   目标二: 摧毁GDI基地=   Objective Two: Destroy the ICBMs targeted at the Philidephia.2   目标二: 摧毁瞄准费城的洲际弹道导弹K   Objective Two: Escort the toxin trucks past the GDI checkpoint to the east.5   目标二: 护送毒素卡车通过GDI检查站向东*   Objective Two: Evacuate the Chameleon Spy.    目标二: 撤离变色龙间谍$   Objective Two: Evacuate the mutants.   目标二: 撤离变种人�   Objective Two: Now find the Mutant Headquarters and knock on their door (attack it!). This should convince Tratos to be sympathetic to our cause.|   目标二: 现在找到变种人总部并敲他们的门（攻击它!）.这应该能说服特拉托斯同情我们的事业*   Objective Two: Remove the GDI trespassers.   目的二: 清除GDI侵入物1   Objective Two: Retrieve the cargo from the train.#   目标二: 从火车上取回货物B   Objective Two: To get production online build a Tiberium Refinery.7   目标二: 建设提矿精炼厂, 实现生产线上化B   Objective Two: Use Toxin Soldiers to "convince" McNeil to join us.=   目标二: 利用毒素步兵"说服"麦克尼尔加入我们   Objective one complete.   目标一完成*   Objective one: Destroy all Nod structures.    目标一: 摧毁所有Nod建筑9   Objective one: Destroy all chemical missile launch sites.,   目标一: 摧毁所有化学导弹发射场.   Objective one: Destroy all the chemical tanks.    目标一: 摧毁所有毒素罐5   Objective one: Remove all Nod presence from the area./   目标一: 清除该区域内的所有Nod势力P   Objective one: Spy on GDI comm center to learn the location of the weapons test.:   目的一: 潜入GDI通信中心, 获取试验场的位置   Objective two complete.   目标二已完成&   Objective two: Capture Vega's Pyramid.#   目标二: 占领维加的金字塔<   Objective two: Capture the train station. DO NOT DESTROY IT!+   目标二: 占领火车站.不要毁了它!5   Objective two: Destroy the Mammoth Mark II prototype.&   目标二: 摧毁猛犸机甲原型机$   Objective two: Destroy the Nod base.   目标二: 摧毁Nod基地V   Once the life form has snacked on the civilian pawns it will feast on the settlements.V   一旦生命体在平民的典当上吃了零食, 它就会在定居点上大快朵颐   Priest: Blessed are the beasts!   牧师: 野兽们有福了!    Priest: Kill the MUTANT invader!'   牧师: 杀了那个顽固的入侵者!   Priest: Kill the Mutant!   牧师: 杀死变种人!9   Priest: Mortimer predicted the coming of these creatures./   牧师: 摩梯末预言了这些生物的到来   Priest: Praise this plant!   牧师: 赞美这棵植物!   Priest: STOP! THIEF!   牧师: 站住! 小偷!   REFINERIES, and SILOS.   炼油厂和筒仓4   Repair the bridge to gain access to the Genesis Pit.    5   Rescue the plebes then take care of those harvesters.)   营救平民, 然后照顾那些收割者   Riot leader neutralized.   暴乱领导人被制服V   Second Objective: "Persuade" the civilians to assist our goal with the Toxin Soldiers.D   目标二: “说服”平民用毒素步兵协助我们实现目标U   Second Objective: Deactivate the firestorm defenses and neutralize the sensor arrays.A   目标二: 关闭火风暴防御系统并使传感器阵列失效'   Second Objective: Destroy CABAL's base.   目标二: 摧毁CABAL的基地6   Second Objective: Destroy the cyborg production plant.&   目标二: 摧毁生化人生产工厂:   Second Objective: Determine if the Kodiak can be salvaged.2   目标二: 确定科迪亚克号是否可以打捞6   Second Objective: Get Dr. Boudreau to the landing pad.+   目标二: 把Boudreau医生送到着陆台E   Second Objective: Maintain ALL factories until reinforcements arrive.5   目标二: 维持所有工厂运作直到援军到达A   Second Objective: Protect food and water processors at all costs.8   目标二: 不惜一切代价保护食品和水加工商#   Second Objective: Repair the array.   目标二: 修复阵列'   Second Objective: Rescue the CIVILIANS.   目标二: 营救平民K   Second Objective: Retrieve a section of CABAL's core from the storage yard.1   目标二: 从堆场取回CABAL岩芯的一部分H   Second Objective: Return the truck containing the Tacitus to the beacon.5   目标二: 把装有塔西佗的卡车送到信标处�   Solomon: Change of plans - We have verified Vega's presence in the pyramid. CAPTURE the pyramid with Vega alive. DO NOT DESTROY IT!�   所罗门:计划改变了——我们已经证实维加在金字塔里.在维加活着的情况下捕捉金字塔.不要毁了它!1   Stop the cargo truck and retrieve the core piece.   停车并取回核心件'   Stop the patrol from alerting the base!    A   Tacitus recovered and loaded on the truck. Proceed to the beacon.,   塔西佗恢复并装上卡车.前往信标.�   Technicians:  We can shut that fencing down for you, just get us into one of the fence power arrays.  The first one is across the water.x   技术人员: 我们可以帮你关掉栅栏, 只要把我们弄到一个栅栏电源阵列里. 第一个在水的对面S   Thanks! We saw something crash to the east. We also spotted a Nod MCV.  Be careful.Z   感谢! 我们看到东边有东西坠落. 我们还发现了一辆Nod基地车. 小心些Y   The life forms are located in a tiberium accelerated staging area called the Genesis Pit.E   这些生命体位于一个被称为创世坑的泰矿加速集结地,   The orders were clear commander - NO DEATHS!-   命令很明确, 指挥官——没有死亡![   The serum within the tranquilizers they use will make them more accommodating to our plans.H   他们使用的镇静剂中的血清会使他们更适应我们的计划$   Third Objective: Assassinate Tratos.   目标三: 刺杀特拉托斯G   Third Objective: Destroy all GDI and civilian structures in the region.5   目标三: 摧毁该地区的所有GDI和民用建筑+   Third Objective: Destroy all Mutant forces.&   目标三: 摧毁所有变种人部队/   Third Objective: Destroy all of CABAL's forces.%   目标三: 摧毁CABAL的所有部队H   Third Objective: Prevent transportation of the last section of the core.,   目标三: 阻止最后一段核心的运输(   Third Objective: Retreat to the Montauk.   目标三: 撤退到蒙托克<   Third Objective: Return the Tacitus to the drop zone beacon.,   目标三: 将塔西佗返回下降区信标   This can't be good.   这不可能是好事J   To bait the Tiberium life forms, lure them out with the drugged civilians.J   通过激怒泰矿生物, 把他们和被麻醉的平民一起引诱出来R   To gain access to the Genesis Pit repair the bridge to the north of your location.;   要进入创世坑, 请修复您所在位置以北的桥梁,   Too many civilian structures have been lost.   失去了太多的民用建筑*   Too many mutant structures have been lost.!   太多的突变结构已经丢失.   Use the ARCHAEOLOGIST to retrieve the Tacitus.!   使用考古学家检索塔西佗:   Use the Mobile EM-Pulse tanks to stop any mutant vehicles.9   使用移动电磁脉冲坦克阻止所有变种人载具,   Use the Toxin soldiers to capture civilians.   使用毒素步兵抓捕平民>   Use the riot troops to force civilians and mutants to retreat.0   使用防暴部队迫使平民和变种人撤退:   Use the truck to transport the Tacitus when you locate it.#   找到塔西佗后, 用卡车运输A   Use your ENGINEER to steal an EVA unit from GDI's RADAR FACILITY.?   让你的工程师从GDI的雷达设施里窃取一个EVA单位%   Villager: My God! Men arm yourselves!'   村民:我的天啊!男人武装自己!)   Villager: Thanks for the warning.  Here's"   村民: 谢谢你的提醒. 这是*   Warning: Do not kill civilians or mutants!'   警告: 不要伤害平民或变种人!C   Warning: Prevent the destruction of mutant and civilian structures.+   警告:防止破坏变种人和民用建筑'   Welcome stranger! Surely the divine one    "   Women and children to the shelter!   妇女和儿童到避难所去!   Zealot: Existance is futile!   狂热者: 存在是徒劳的!   Zealot: I'm coming to join you!   狂热者:我来加入你们!   Zealot: Kill the Heretics!   狂热者: 杀了异教徒!   Zealot: Look! A Mutant!   狂热者:看!变种人!3   Zealot: Mutant Abomination! How dare you defile the,   狂热者:变种人灭绝!你怎么敢玷污(   Zealot: Wha?! They've killed the Leader!$   狂热者: 什?! 他们杀了首领!   a reward for your concern.   感谢你的关心)   actively capturing civilians to turn them   积极抓捕平民+   all dead.  Concentrate on those harvesters.)   都死了. 集中精力对付那些矿车"   and an MCV will be sent in to you.   CABAL: 届时将派遣MCV支援*   currently harvesting biological components   目前正在收获生物成分	   en route.   途中(   evacuate the city immediately!  CABAL is   立即撤离城市! CABAL是(   everyone is evacuated.  Please take this(   所有人都被撤离了.请收下这个    for his Cyborgs. Arm Yourselves!#   为了他的机器人.武装自己!,   has guided your footsteps to this Holy Land.$   指引你的脚步来到这片圣地   humans into his Cyborg army.$   人类加入了他的赛博格军队!   humans to turn them into Cyborgs.   把人类变成变种人   into Cyborgs.   进入Cyborgs.   is so pleased that they have consented to send   很高兴他们同意发送,   off now.  Extraction in T minus two minutes.    *   operations in this sector and is capturing!   该领域的业务正在被占领%   rejoice in the glory of our savior...'   为我们救世主的荣耀欢舞吧...   sanctity of our Holy ground?   我们圣地的神圣性?   storm abates.   暴风雨减弱了/   that we aid these Civilians.  We cannot refuse.        the JUGGERNAUT. Do not waste it.   神像.不要浪费它   to help in your battle.   来帮助你战斗$   will alert Hassan to their presence.   会提醒哈桑他们的存在
   you a MCV.   你一个基地车   you more funding.   你有更多的资金strings    �  :     -DESTNET = Specify Network Number of destination system
+    -DESTNET = 指定目标系统的网络号
5     -MESSAGES = Allow messages from outside this game.
/    -MESSAGES = 允许来自游戏外部的消息
*     -SOCKET = Network Socket ID (0 - 16383)
(    -SOCKET = 网络 Socket ID (0 - 16383)
2     -STEALTH = Hide multiplayer names ("Boss mode")
3    -STEALTH = 隐藏多人游戏名称("Boss模式")

   %d Credits   %d 分   %d Starting Units   %d 启动单位   %s
%s
Rank : %d   %s
%s
排名 : %d   %s
Rank : %d   %s
排名 : %d   %s Accessibility   %s 可访问性	   %s Cities	   %s 城市	   %s Cliffs	   %s 悬崖   %s Hills	   %s 山丘   %s Tiberium	   %s 泰矿   %s Tiberium Fields   %s 泰矿田   %s Vegetation	   %s 植被   %s Water	   %s 水体   %s changed game options!   %s 改变了游戏选项!   %s declares war on %s   %s 向 %s 宣战!   %s has allied with %s   %s 与 %s 结盟!#   %s has been banned from the channel   %s 已被禁止进入该频道!   %s has been defeated!   %s 被击败了!   %s has formed a new game.   %s 开了一个新游戏   %s has left the game.   %s 离开了游戏   %s playing %s   %s 正在游戏 %s%   %s proposes kicking %s from the game.   %s 建议将 %s 踢出游戏	   %s's Game   %s 的游戏   %s's game is now in progress.   %s 的游戏正在进行中   (NOT USED ANYMORE)   (不再使用)
   -- More --
   --更多--  A cyborg commando has been sent to retrieve you.  Once free, rendezvous with your rescue team to the south.  Use them to locate and free Oxanna before she is transported to the main GDI facility.  After she has been freed, capture a GDI transport to make your escape.  �   一个生化尖兵被派去营救你, 逃出之后尽快在南边集合. 在奥克斯安娜被转移到GDI的主要设施之前, 尽快解救她. 解救她后, 拦截一辆GDI运输车用于撤离.-   A mouse is required for playing Tiberian Sun.1   游玩《泰伯利亚之日》需要一只鼠标.(   A required field is missing, or invalid.   必填字段缺失或无效.�   A sensor net protects the valley where Tratos is being held.  To facilitate his rescue, we must disable the array that controls this highly sensitive net.  Once down, it will be much easier to get Tratos out of the valley.�   一片传感器网络保护着特拉托斯被关押的山谷. 为了便于营救他, 我们必须关闭这个网络的控制阵列, 这样再把特拉托斯带出山谷会容易得多.   Abundant	   丰富的   Abundant Tiberium   丰富的泰矿   Abundant Water   丰富的水   Accepted	   已接收	   Activated	   已激活   Add Select Team %2d   添加选择队伍 %2d	   Afternoon   下午   All Locations   所有位置0   All users must accept before the game can start..   所有玩家必须都接受才能开始游戏.   Alliance   联盟)  An upgrade is required for this game
Do you want to download it now?
 
 
Warning: use of "trainers", third-party cheat programs, or any other modification of Tiberian Sun may cause the automatic update procedure to fail. Please remove any such programs or reinstall Tiberian Sun before continuing.	  游戏当前需要升级
你想立即下载吗?


警告: 使用"trainers"第三方作弊程序, 或任何其他修改泰伯利亚之日的程序都可能会导致自动更新失败. 请在继续之前删除任何此类程序或重新安装《泰伯利亚之日》.#   Analyzing combat zone topography...   分析战区地形...�  Another possible location of the fighter production facility.  Use the mutants to locate the position of the fighter production facility.  They must remain undetected. If Nod suspects enemy forces, they will cloak their production facility and deploy troops.  If the mutants can hide from the Nod troops for a short period, Nod will assume the area is clear, and uncloak the base.  Once we have recorded the location of the base, the mission will be complete.+  战斗机生产设施的另一个可能位置. 利用变种人确定该设施的位置, 他们必须保持隐蔽. 如果Nod起疑, 他们会使设施隐形并部署部队, 尽量让变种人及时躲避Nod部队, 以避免惊扰他们. 只要我们记录了该设施的位置, 任务就算完成了.   Answering Canceled   应答已取消   Answering...   正在应答...   April   四月>   Are you sure you want to remove user '%s' from the login list?2   您确定要从登录列表中删除用户"%s"吗?6   Are you sure you want to reset the hotkey assignments?%   您确定要重置快捷键分配吗?	   Atom Bomb	   原子弹   August   八月   Back   返回   Bad   坏的
   BattleClan
   BattleClan   BattleClan Game   BattleClan 游戏�   Be advised, the Brotherhood will attempt to destroy the impact site.  GDI reinforcements are en route.  Protect the site until they arrive.j   注意, 兄弟会将试图摧毁坠机现场. GDI增援部队正在赶来, 保护现场直到他们到达.�   Be advised: Kane is determined to destroy you.  The ion storm has grounded the Kodiak.  We must protect it until the storm abates.  Production will be limited.  There is a high probability of equipment malfunction.  Caution is advised.�   注意: 凯恩已下决心要消灭你. 离子风暴使科迪亚克停飞, 我们必须保护它直到风暴减弱. 你的生产将受到限制, 设备故障的可能性很高, 建议谨慎行事.   Best Scores   最佳成绩   Blue   蓝色   Bridges Destroyable   可摧毁桥梁	   Buildings   建筑   Bytes read: %d / %d.   字节读取: %d / %d.-   Bytes read: %d / %d.    Time left: %d seconds+   字节读取: %d / %d.  剩余时间: %d秒
   CASUALTIES   伤亡   CURRENCY   资金   CUSTOM -   自定义 -   Cancel   取消   Center Base   居中基地   Center Team %2d   居中队伍 %2d   Center View   居中视图1   Center the tactical view on the last radar event.4   把战术视野居中在最后一次雷达事件上.)   Center the view about selected object(s).   将选定对象的视图居中.(   Center the view about the player's base.%   将玩家基地周围的视图居中.   Channel Operator   频道运营商   Charging...   填充中...   Chat Server Error   聊天服务器错误R   Check your connection to the internet.  If you were disconnected from the internet>   检查你的互联网连接. 如果你与互联网断开连接   Civilian Building   民用建筑8   Click cancel to abort this game and return to the lobby.-   单击"取消"中止此游戏并返回大厅.>   Click on a name to propose removing that player from the game.<   点击一个名字, 以提出将该玩家从游戏中删除.   Click to Continue   点击继续(   Compensating for ambient light values...   环境光补偿值...    Compiling wartime conventions...   编纂战时公约...�   Complete destruction of the missile complex is essential.  Be advised, Nod will use their Tiberium missiles and their new fighter prototypes against you.q   彻底摧毁导弹设施至关重要. 请注意, Nod将使用他们的泰矿导弹和原型战斗机来对付你.   Computer   电脑   Connecting to Westwood Online   连接到Westwood网络   Connecting...	   连接...?   Connection error! Check your cables. Attempting to Reconnect...7   连接错误! 请检查网线. 并尝试重新连接...   Connection error! Redialing...   连接错误! 重新拨号...%   Connection error! Waiting for Call...   连接错误! 等待来电...?   Connection to %s has been interrupted. Attempting to reconnect.0   与 %s 的连接已中断. 尝试重新连接...   Connection to %s lost!   与 %s 的连接丢失!   Continue   继续   Control   控制:  Control of the mutants is in our grasp.  Their headquarters is located to the north of your drop-off position.  The GDI units you will need to implicate in this deception occupy a small base to the southwest.  Do not mar the Brotherhood's name any further.  Allow the blame to fall squarely on Solomon's shoulders.�   我们已经控制了变种人, 他们的总部在你下车位置的北面. 而你要诱骗的GDI部队占据了西南部的一个小基地. 不要再玷污兄弟会的名声了, 就让所罗门来承担这些吧.E   Could not connect to Westwood Online, check your Internet connection.;   无法连接到Westwood网络, 请检查您的网络连接.V   Could not connect to the World Domination Tour server, or there is no server availableJ   无法连接到世界统治之旅服务器, 或者没有可用的服务器   Could not create the channel   无法创建频道   Couldn't get the server list   无法获取服务器列表   Couldn't page user   无法分页用户   Create Team %2d   创建队伍 %2d   Created channel: %s   已创建频道: %s.   Creates Team %d from currently selected units.'   从当前选定的单位创建团队%d.)   Creating theories on likely enemy plan...!   对可能的敌人设定计划...   Credits:   资金:   Cyan   青色   Data Queue Overflow   数据队列溢出   Day : %d   天: %d   December	   十二月   Default   默认   Delete Waypoint   删除路径点   Delete selected waypoint.   删除选定的路径点.   Delete this file?   删除此文件?   Deploy Object   部署对象   Deploy selected object(s).   部署所选对象."   Deploying forces to combat zone...   向战区部署部队...   Desert   沙漠%   Destination game version is outdated.   目标游戏版本已过时.=   Destination network address must be in the format xx.xx.xx.xx/   目标网络地址的格式必须为xx.xx.xx.xx   Destroy all enemy units   摧毁所有敌方单位   Destroy all enemy units.   摧毁所有敌方单位.�   Destroying the base in this sector will prevent further removal of artifacts from the crash site.  In addition, Nod will not be able to reinforce the site from this location.�   摧毁该区域的基地将阻止Nod进一步从坠机现场搬运外星遗物. 同时, Nod也将无法从此地向外派遣增援._   Destroying the supply base here will prevent the missile complex from receiving reinforcements.@   摧毁这里的补给基地可以阻止导弹基地得到增援.   Dialing Canceled   拨号已取消
   Dialing...   正在拨号...   Display game options dialog.   显示游戏选项对话框.   Downloading file %d of %d...   正在下载文件 %d 的 %d...   Dusk   黄昏   EM Pulse   电磁脉冲   Easy   简单   Economy   经济   Enemy Soldier   敌方步兵   Enemy Structure   敌方建筑
   Enemy Unit   敌方单位G  Enter the sector and deploy your base.  Once you have established a tiberium waste facility, convoys of tiberium waste will begin arriving.  Protect the convoys at all cost.  Once we have enough tiberium waste, the missile will be ready for use against GDI.  Destroying their base, once it is infected, will be a simple matter./  进入区域并部署您的基地. 当你建立了泰矿回收厂之后, 一支泰矿回收车队就会开始出发. 不惜一切代价保护这支车队. 只要我们有了足够的泰矿, 就可以用来制造导弹对付GDI. 一旦他们的基地被污染, 摧毁它将是一件极其简单的事情.7   Error - Modem did not respond to initialisation string.7   错误 - 调制解调器没有响应初始化字符串.l   Error - Modem failed to respond to compression disable command. Your Windows configuration may be incorrect.[   错误 - 调制解调器未能响应压缩禁用命令. 您的Windows配置可能不正确.j   Error - Modem failed to respond to compression enable command. Your Windows configuration may be incorect.[   错误 - 调制解调器无法响应压缩启用命令. 您的Windows配置可能不正确.q   Error - Modem failed to respond to error correction disable command. Your Windows configuration may be incorrect.a   错误 - 调制解调器未能响应错误纠正禁用命令. 您的Windows配置可能不正确.p   Error - Modem failed to respond to error correction enable command. Your Windows configuration may be incorrect.[   错误 - 调制解调器未能响应纠错启用命令. 您的Windows配置可能不正确.e   Error - Modem failed to respond to flow control command. Your Windows configuration may be incorrect.X   错误 - 调制解调器未能响应流控制命令. 您的Windows配置可能不正确.$   Error - Modem returned error status."   调制解调器返回错误状态.%   Error - TIme out waiting for connect.   错误 - 等待连接超时.6   Error - Too many errors initialising modem - Aborting.:   错误 - 初始化调制解调器时错误太多 - 中止.,   Error - Unable to disable modem auto answer.1   错误 - 无法禁用调制解调器自动应答.%   Error - Unable to set the video mode."   错误 - 无法设置显示模式.;   Error - other player does not have this expansion scenario..   错误 - 其他玩家没有这个扩展场景.   Error in the InitString   初始化字符串错误   Error joining channel %X   加入频道 %X 出错   Error loading game!   加载游戏时出错!   Error saving mission!   保存任务时出错!'   Failed to initialize. Please reinstall.!   初始化失败, 请重新安装.   Fast   快   Faster   更快   Fastest   最快   February   二月*   Fetching World Domination Tour information   获取世界统治之旅信息   Fetching ladder information   获取梯子信息   Fetching server list   正在获取服务器列表   Fetching squad information   获取小队信息   Few   少
   Few Cities   少量城市
   Few Cliffs   少量悬崖	   Few Hills   几座小山   Few Tiberium Fields   少量泰矿   Final analysis of outcome...   结果的最终分析...   Find failed   查找失败   Finding Patch...   寻找补丁...	   Firestorm   火焰风暴   Firestorm BattleClans   火焰风暴BattleClans   Firestorm Defense Toggle   火焰风暴防御开关   Firestorm Players   火焰风暴玩家,   Firestorm must be enabled to join this game..   必须启用火焰风暴才能加入此游戏.%   Firestorm required to join this game.%   加入这个游戏需要火焰风暴.
   Fog of War   战争迷雾   Follow   跟随   Four Player Only   仅限四人(   From Computer: It's just you and me now!'   来自电脑: 现在只有你和我了!   GDI Barracks	   GDI兵营   GDI Comm. Center   GDI通信中心   GDI Tech Center   GDI 科技中心	   Game Over   游戏结束了   Game has a password   游戏有密码   Game is closed.   游戏已关闭.   Game is full.   已经满员了.\   Game versions incompatible. To make sure you have the latest version, visit www.westwood.comP   游戏版本不兼容. 为确保您拥有最新版本, 请访问www.westwood.com   Game was cancelled.   游戏被取消了   Game# %d   游戏#  %d   Game: %d
   游戏: %d'   Gathering intel on involved factions...   收集相关派系的情报...   Gold   金色   Goodie Crates   物资板条箱   Goto Radar Event   跳转雷达事件   Gray   灰色   Green   绿色   Guard	   警戒的   Hand of NOD	   NOD之手   Hard   困难   Harvester Truce   采矿车休战@  Hassan communicates to the Brotherhood through a nearby TV station.  With the Brotherhood in chaos, the opportunity to divide Hassan from his followers presents itself.  Capture the TV station and those once loyal to Kane's technology of peace will return to the fold.  And as for Hassan's pathetic guards -- crush them.  哈桑通过附近的电视台与兄弟会联系. 随着兄弟会陷入混乱, 哈桑与追随者之间也出现了隔阂. 占领电视台, 这样那些曾经热衷于凯恩科技的人就会重返正轨. 至于哈桑那些可怜的守卫... 把他们干掉!   Heavy   重   Heavy Vegetation   厚重的植被   High   高   High Accessibility   高可访问性
   Host Rank:   房主排名:   Huge Map	   大地图   IPX not available   IPX不可用   IRQ already in use   IRQ已在使用中Q   If all other players have connection times in the red then you have probably beenY   如果所有其他玩家的连接时间都是红色的, 那么有问题的很可能是你   Ignore   忽略   Ignore User   忽略用户�   Impulse signatures emanating from Cairo suggest Kane will launch his world-altering missile within hours.  You must destroy the pyramid temple before he has the chance to launch.  There are no alternatives.�   来自开罗的脉冲信号表明, 凯恩将在数小时内发射足以颠覆世界的导弹. 你必须在他发射导弹之前摧毁金字塔神殿, 我们别无选择.�   In this sector lies a Nod base overrun with tiberium-based lifeforms.  Find the base, reactivate it, and use the tiberium life to fill our missiles.  When you have enough of the tiberium substance, launch the missile against the GDI base and destroy it.�   在这个区域, 有一个泰伯生命体泛滥的Nod基地. 找到基地并重新激活它, 用泰伯生命体充能我们的导弹. 当你有足够的泰矿物质时, 向GDI基地发射导弹并摧毁它.A   Incompatable scenario file detected. The scenario may be corrupt.9   检测到不兼容的场景文件. 场景可能已损坏.   Indestructable Bridges   不可摧毁的桥梁   Infantry   步兵   Initializing Modem...Standby!   初始化调制解调器...就绪w   Insufficient disk space to save a game.  Please delete a previous saved games to free up some disk space and try again.h   磁盘空间不足, 无法保存游戏. 请删除以前保存的游戏释放一些磁盘空间后再试.	   Interface   界面   Invalid Port or Port is in use$   端口无效或端口正在使用中(   Invalid Port/Address. COM 1-4 OR ADDRESS   COM端口1-4或地址无效.   Invalid option switch.   无效的选项开关.   Invalid/Missing   无效/缺失
   Ion Cannon	   离子炮�   It is highly probable that the Brotherhood will attempt to remove technology from the crash site and store it at the technology center.  Locate and secure the crash site, then capture the technology center.�   兄弟会极有可能试图从坠机现场提取技术并将其存储在技术中心. 找到并保护坠机现场, 然后占领Nod技术中心.�  It is imperative that you prevent the train from reaching the Nod base.  Remember, destroying the locomotive will immediately stop the train.  Recent ice melts in the region have disabled the only train bridge.  You must move quickly as Nod engineers are on their way to repair it.  The crystals can be recovered easily if you get to the train before Nod can repair the bridge.  Otherwise, we will need to attack the base in order to reclaim the crystals.E  你必须阻止火车到达Nod基地. 记住, 摧毁火车头会使火车立即停止. 该地区融化的冰瘫痪了唯一的火车桥. 你必须快速行动, 因为Nod的工程师正在修理它的路上. 如果你在Nod修好桥之前到达火车, 就能轻松抢走水晶. 否则, 我们就得进攻Nod基地夺回水晶.   January   一月   Join   加入   Joining Lobby   加入大厅   Joining channel: %s   加入频道: %s   July   七月   June   六月�  Kane's vision is at hand.  Unfortunately GDI's orbital station, the Philadelphia, can stop the missile that will take us into the future.   We must destroy the Philadelphia at all costs!  The Philadelphia will require three orbits over this sector before it can locate our missile.  You must get three ICBM launchers into position before the Philadelphia's final orbit is complete.  With the ICBMs in place, we can bring GDI's command station down.  All this remains contingent, of course, on McNeil's helpfulness.  You must pretend to pursue him back towards the GDI base.  They will open the perimeter to let him in.  Once he is in, he will deactivate the perimeter shortly thereafter.  凯恩的愿景就在眼前了. 不幸的是, GDI的费城空间站可以拦截我们的导弹. 我们必须不惜一切代价摧毁空间站! 这座空间站需要在这个区域上空飞行至少三圈, 而在空间站到达最终轨道之前, 你必须将三个导弹发射器就位. 有了洲际弹道导弹, 我们就可以摧毁GDI的指挥中心. 当然, 这一切都取决于麦克尼尔的配合. 你需要假装追击他, 促使GDI让他进入基地. 一旦他成功潜入, 很快就会打开大门放我们进去.   Kills   杀死击杀   Kills:   击杀:   Large   大	   Large Map	   大地图   Leave   离开
   Line busy.   线路繁忙.   Lobby   大厅   Logging off Westwood Online   注销Westwood网络   Losses   损失O   Lost connection to Westwood Online, outside users will not be able to page you.B   与Westwood Online的连接中断, 外部用户将无法呼叫您.   Low   低   Low Accessibility   低可访问性	   Low Power   电力不足   MCV Not Redeployable   MCV不可重新部署   MISSION EFFICIENCY   任务效率   MISSION TIME LAPSE   任务用时   Many   许多   Many Cities   许多城市   Many Cliffs   许多悬崖
   Many Hills   许多山丘   Many Tiberium Fields   许多泰矿
   Map Error!   地图错误!   Map: %s
   地图: %s   March   三月   May   五月   Medium   中   Message:   消息:   Mission Accomplished   任务已完成   Mission Failed   任务失败   Mission Saved   任务已保存"   Mission is loading. Please wait...   正在加载任务.请稍等...   Mission saving - Please Wait...   任务保存中 - 请稍等...   Mode   模式   Morning   早晨   Multi-Engineers   多位工程师   Multiplayer Game   多人游戏   Mutated	   突变的   NOD Barracks	   NOD兵营   Name:   名称:
   Narrow Map   缩小地图   New   新建   New Chat	   新聊天   New Game	   新游戏   Next Object   下一个对象   Night   夜晚   No   否   No Goodie Crates   没有物资板条箱   No Sound Card Detected   没有检测到声卡   No Starting Bases   无起始基地   No carrier.
   无载波.M   No dial tone. Ensure your modem is connected to the phone line and try again.P   没有拨号音. 确保调制解调器已连接到电话线, 然后再试一次.   No preview available.   没有可用的预览.�  Nod has taken over much of our Hammerfest base in their search for the disrupter. Nod has reactivated the perimeter to prevent GDI from attacking.  Water assault remains your only option.  Find the Firestorm Defense structure generating the perimeter and deactivate it.  Only then can reinforcements arrive.  Proceed to destroy Nod's primary base, and prevent them from attacking again.D  Nod为了寻找声波坦克, 夺取了我们哈默菲斯特基地的大部分. Nod已经重新激活了防线, 以防止GDI攻击. 从水上进攻仍然是你唯一的选择, 找到周边的"火焰风暴"防御建筑并将其关闭. 只有这样, 增援部队才能到达. 摧毁Nod的主要基地, 防止他们再次进攻.   Normal   正常   Normal Engineers   普通工程师A   Not a Null Modem Cable Attached! It is a modem or loopback cable.N   没有一个调制解调器电缆连接! 它是调制解调器或环回电缆.   Nothing to join!   没什么可加入!   November	   十一月   Number invalid.   号码无效.   Numerous Cities   许多城市   Numerous Cliffs   大量悬崖   Numerous Hills   许多山丘   Numerous Tiberium Fields   大量泰矿   OK   确定   October   十月   Off   关   Official chat channels   官方聊天频道   On   开   On Hold   等待j  One of two possible locations for the fighter production facility.  Use the mutants to locate its whereabouts while remaining undetected.  If detected, Nod will cloak the factory and deploy more troops.  Hide the mutants, and Nod will once again uncloak their base.  After the base location is recorded, GDI dropships will immediately arrive with reinforcements.  战斗机工厂有两个可能的地点. 利用变种人定位它的位置, 同时不被发现. 如果被发现, Nod将隐藏工厂并部署更多部队, 此时隐蔽变种人, 等待Nod暴露工厂. 在工厂位置被记录下来后, GDI运输船将立即带着增援部队抵达.@   One or more DLL files were missing
or damaged. Please reinstall.9   一个或多个DLL文件丢失或损坏.
请重新安装.   Only one player?   只有一个玩家?%   Only the host can modify this option."   只有房主可以修改此选项.   Oops!   哦欧!   Options   选项   Options Menu   选项菜单   Orange   橙色   Other game channels   其他游戏频道   Other system not responding!   其他系统没有响应!   Overwrite existing save game?   覆盖已保存的游戏?   Packet received too late!   收到数据包太晚了!	   Page User    1   Page a Westwood Online user. (Internet play only)8   为Westwood网络用户添加页面.(仅限网络游戏)%   Page sidebar selection list downward.   侧边栏选择列表向下.#   Page sidebar selection list upward.   侧边栏选择列表向上./   Page sidebar structure selection list downward."   页面侧边栏建筑列表向下.-   Page sidebar structure selection list upward."   页面侧边栏建筑列表向上.*   Page sidebar unit selection list downward."   页面侧边栏单位列表向下.(   Page sidebar unit selection list upward."   页面侧边栏单位列表向上.   Page was successful.       Parameters:
   参数:
   Pink   粉色3   Player %s has changed the connection speed setting.&   玩家 % s已更改连接速度设置.-   Player %s has changed the game speed setting.    玩家 %s 已更改游戏速度.   Players   玩家   Please Choose Map   请选择地图   Please Stand By...   请稍候...   Please enter a message to send   请输入要发送的消息/   Please insert CD %d (%s) into the CD-ROM drive.%   请将CD %d(%s)插入CD-ROM驱动器.6   Please insert a Tiberian Sun CD into the CD-ROM drive.@   请在CD-ROM驱动器中插入《泰伯利亚之日》的光盘.7   Please select 'Settings' to setup default configuration&   请选择"设置"以还原默认配置   Poor   贫瘠   Power = %d
Drain = %d   电力 = %d
负载 = %d
   Power Mode   电源模式   Previous Object   上一个对象   Pri.   主.   Primary   主要   Proceeding with audio disabled.   关闭音频继续.   Purple   紫色   Radar Toggle   雷达开关
   Random Map   随机地图   Rank   排名   Ready   就绪   Receiving scenario from host.   从主机接收场景.   Reconnection Error!   重连错误!   Red   红色   Redeployable MCV   可重新部署MCV   Reject   拒绝   Release   释放   Repair Mode   修复模式   Request denied.   请求被拒绝.   Requesting channel list   请求频道列表   Requesting new login...   正在请求新登录...   Resume Mission   恢复任务   Reviewing History
   回顾历史
   SEARCHING...   正在搜索...   Scarce   稀缺   Scarce Tiberium   稀缺的泰矿   Scarce Water   稀缺的水   Scatter   分散   Scatter selected object(s).   分散选定对象.	   Scenario:   场景:   Scenarios don't match.   场景不匹配   Score   得分   Screen Capture   截屏   Scroll East   向东滚动   Scroll North   向北滚动   Scroll South   向北滚动   Scroll West   向西滚动'   Scroll sidebar selection list downward.   向下滚动侧边栏列表.1   Scroll sidebar structure selection list downward."   向下滚动侧边栏建筑列表./   Scroll sidebar structure selection list upward."   向上滚动侧边栏建筑列表.,   Scroll sidebar unit selection list downward."   向下滚动侧边栏单位列表.*   Scroll sidebar unit selection list upward."   向上滚动侧边栏单元列表.    Scroll tactical map to the east.   向东滚动战术地图.!   Scroll tactical map to the north.   向北滚动战术地图.!   Scroll tactical map to the south.   向南滚动战术地图.    Scroll tactical map to the west.   向西滚动战术地图.&   Scrolls sidebar selection list upward."   向上滚动侧边栏选择列表.   Searching for %s....   正在搜索 %s ....!   Secondary check of combat zone...   作战区域二次检查...   Select Same Type   选择相同类型   Select Team %2d   选择队伍 %2d   Select View   选择视图-   Select all owned objects in the current view.+   选择当前视图中所有拥有的对象.%   Select and center view about team %d.   选择并居中查看队伍 %d.:   Select members of team %d without unselecting other units.:   选择队伍 %d 的成员, 而不取消选择其他单位.   Select members of team %d.   选择团队 %d 的成员.   Select the next object.   选择下一个对象.   Select the previous object.   选择上一个对象.	   Selection   选择9   Selects all units of the same type as currently selected.1   选择与当前所选类型相同的所有单位.	   Sell Mode   出售模式*   Sending GO acknowlegement - Please Wait...#   正在发送GO确认 - 请稍候...#   Sending GO request - Please Wait...   发送GO请求 - 请等待...#   Sending scenario to remote players.   向远程玩家发送场景.	   September   九月   Set Bookmark 1   设置书签 1   Set Bookmark 2   设置书签 2   Set Bookmark 3   设置书签 3   Set Bookmark 4   设置书签 42   Set the selected object(s) into 'guard area' mode.*   将所选对象设置为"保护区"模式.!   Set view bookmark map position 1.!   设置视图书签地图位置 1.!   Set view bookmark map position 2.!   设置视图书签地图位置 2.!   Set view bookmark map position 3.!   设置视图书签地图位置3 .!   Set view bookmark map position 4.!   设置视图书签地图位置 4.   Settings   设置   Short & Wide Map   短宽地图
   Short Game   快速游戏	   Short Map	   短地图   Sidebar	   侧边栏   Sidebar Down   侧边栏向下   Sidebar PageDown   侧边栏向下翻页   Sidebar PageUp   侧边栏向上翻页
   Sidebar Up   侧边栏向上   Signing off - Please Wait...   结束广播 - 请稍候...�   Since you are under the age of 13 our privacy policy requires that you send us a parental consent form to continue.  Press 'yes' to open your web browser to this page.u   由于您未满13岁, 我们的隐私政策要求您发送家长同意书才能继续. 点击"是"以打开浏览器.   Sky Blue	   天蓝色   Slow   慢   Slower   更慢   Slowest   最慢   Small   小	   Small Map	   小地图)   Socket number must be between 0 and 16383*   套接字号码必须介于0和16383之间0   Sorry, that player or rank is not in the ladder.0   对不起, 那个玩家或级别不在天梯上.   Sparse   稀疏   Sparse Vegetation   稀疏的植被   Spy Info   间谍消息   Starting Bases   起始基地   Stop   停止   Stop Object   停止对象   Stop the selected object(s).   停止所选对象.   Structure List Down   建筑列表向下   Structure List PageDown   建筑列表向下翻页   Structure List PageUp   建筑列表向上翻页   Structure List up   建筑列表向上
   Structures   建筑	   Surrender   投降   Taiga	   针叶林a   Take a snapshot of the game screen. (Saved as 'SCRNxxxx.PCX' file in Tiberian Sun run directory.)\   拍摄游戏屏幕的快照 .(另存为泰伯利亚之日目录中的"SCRNxxxxx.PCX"文件.)�   Taking out this weak GDI position will allow us to reclaim our Sarajevo temple without interruption.  Move in under the cover of an ion storm when GDI's communications will be down.  Take out the comm center before the storm subsides.�   消灭这个脆弱的GDI据点将使我们能够不受干扰地夺回我们的萨拉热窝神殿. 趁GDI通讯中断时, 在离子风暴的掩护下行动. 在风暴平息前摧毁通讯中心.�   Taking out this weak GDI position will allow us to reclaim our Sarajevo temple without interruption.  Move to an open area and build your base.  GDI patrols are known to be in the area.  Do not mar the brotherhood's name any further.�   消灭这个脆弱的GDI据点将使我们能够不受干扰地夺回我们的萨拉热窝神殿. 前往开阔的地方建立你的基地. 已知GDI巡逻队在该地区, 不要再玷污兄弟会的荣耀了.   Tall & Narrow Map   高窄地图   Tan       Team   队伍   Tech Level %d   科技等级 %d
   Technician	   技术员	   Temperate	   温和的   Temple of NOD
   NOD 神殿   That channel is full   那个频道已经满了   That game channel has closed!   那个游戏频道已经关闭了!   That login is already being used.   该登录已被使用.%   That login or password was incorrect.   该登录名或密码不正确.�  The GDI defense perimeter is located here.  Do not destroy any GDI factories during your assault - you will need them to build GDI units under our control.  Once Jake McNeil's inspection detail is in our converted base, attack!  Kill all but McNeil.  Use the special toxin soldiers provided to control McNeil.  Once he has been "persuaded" to help us in our cause, EVAC him as directed.  If he detects the trap, capture him before he can flee the sector.   �  GDI哨所位于这里, 你在进攻时不要摧毁任何GDI工厂 - 你需要利用它们建造GDI的单位. 一旦确认杰克·麦克尼尔到达被我们改建的基地, 就发动攻击! 杀了除麦克尼尔的所有人. 使用特殊的毒素步兵来控制麦克尼尔, 当他被"说服"加入我们的事业后, 就按照计划撤离他, 如果他发现这是陷阱, 那就在他逃跑之前抓住他.H  The Nod forces that attacked our Phoenix base are in this sector.  Their base must be destroyed in order to secure the region.  However, there is a significant civilian population requiring evacuation.  GDI transports will evacuate the civilians once all Nod SAM sites are destroyed.  The Nod base can then be safely terminated.  袭击费城基地的Nod部队就在这个区域. 他们的基地必须被摧毁, 以确保该地区的安全. 但是, 有大量平民需要撤离. 当所有Nod导弹基地被摧毁后, GDI运输车就会撤离平民, 之后就可以安全地清除Nod基地.   The Westwood online support library is either missing or invalid. Please reinstall the shared internet components from your CD.T   Westwood在线支持库缺失或无效. 请从CD重新安装共享的internet组件.N   The World Domination Tour information was either not downloaded or is corrupt..   世界统治之旅信息未下载或已损坏.[   The active World Domination Tour territories have changed.  Relocating to new front line...P   世界统治之旅的活跃地区已经发生了变化, 搬迁到新的前线...  The alien craft is located in this region - find it!  You must utilize your stealth advantage, as the area is infested with GDI.  Once the craft is located, get an engineer inside to retrieve the Tacitus.  Should you encounter Vega's forces, consider them expendable.�   外星飞船就在这个地区 - 找到它! 你必须利用你的隐形优势, 因为这个地区到处都是GDI. 一旦找到飞船, 派一名工程师进去取回塔西佗. 如果你找到维加的部队, 别怕浪费, 他们是可以牺牲的.&   The channel ban on %s has been removed"   对 %s 的频道禁令已被移除~   The display mode will be changed. If there is a problem with the new display mode then wait and the old mode will be restored.P   显示模式将更改. 如果新显示模式有问题, 请等待恢复旧模式.F   The download failed, please check your connection and try again later.2   下载失败, 请检查您的连接, 稍后重试.@   The host has changed game options, press accept if you're ready.D   房主已更改游戏选项, 如果您准备好了, 请点击接受.   The host has selected   主机已选择b   The infidel Hassan has been tracked to this region of Cairo.  Build a base and remove the usurper.\   异教徒哈桑被追踪到开罗的这个地区. 建立一个基地, 除掉这个篡位者.;  The informant must make contact with the mutants south of the GDI base.  Use the mutants to protect the informant and to eliminate GDI patrols.  Reinforcements will arrive after you have secured the railway tunnel here.  Use them to locate and destroy the research facility.  The mutants, of course, are expendable.�   线人必须与GDI基地以南的变种人取得联系. 利用变种人来保护线人, 并消灭GDI巡逻队. 等你把这里的铁路隧道修好后, 援军就会到达. 用它们来摧毁研究设施. 当然, 变种人也是可以牺牲的.�   The installed version of the Westwood Online support library is too old. Please reinstall the shared internet components from your CD.[   Westwood Online支持库的安装版本太旧. 请从CD重新安装共享的internet组件.�  The large dams that power Vega's base lie in this sector.  Destroying them will temporarily drain power from his base.  To aid you in your objective, attack his island facility before he can bring new generators online.  The dam can be destroyed by disabling the two regulator stations in this sector.  GDI air support will be available if you can find a way to contact them and confirm your target. c  为维加的基地供电的大型水坝就在这个区域. 摧毁它们会暂时中断敌人基地的能源. 为了帮助你完成目标, 在他把新的发电机上线之前攻击他的岛上设施. 大坝可以通过关闭该区域的两个调节站而被摧毁. 如果你能找到与GDI空军联系的方法, 那么你可以得到他们的空中支援.  The mutant female may be trying to reach the underground railway system located in New Detroit.  Move in and control the station before she arrives.  If she boards the train, you must stop it immediately.  This may be our last chance of capturing the abomination.�   这个女变种人可能正试图到达位于新底特律的地下铁路系统, 我们要在她到达之前控制车站. 如果她登上了火车, 你必须立即将其拦截, 这可能是我们抓住这可憎之物的最后机会.^  The mutants are being held on an island in this sector.  We can spare a small force to attempt a rescue.  The area leading to the island is heavily guarded.  If you are detected, more Nod forces will arrive.  Avoiding Nod patrols is advised.  You must rescue all ten mutants and lead them to the dust-off zone.  Periodic airstrikes will be available.=  变种人被关押在这里的一个岛上, 我们可以抽出一小部分力量去营救. 通往该岛的区域戒备森严, 如果你被发现, 更多的Nod部队将会到达. 建议避免与Nod巡逻队接触. 你必须营救所有变种人, 并将他们带到撤离区, 同时我们将定期对敌人进行空袭.%   The requested color is already taken.   请求的颜色已采用.M  The train transporting the mutants is headed to this power grid.  The grid powers the missile complex.  Merely destroying the grid is inadequate: Nod will compensate by building more power plants at the base.  Use all the mutants to plant C4 charges on all the power plants.  We'll detonate the C4 when we attack the missile complex.  运送变种人的火车正驶向这个电网. 这个电网为导弹阵列供电力. 但仅仅摧毁电网是不够的: Nod将通过在基地建造更多的发电厂来弥补. 派遣变种人在所有发电厂上安装C4炸药, 当我们向导弹系统发动攻击时再引爆.;   There are already 2 players with your serial# in that game.8   游戏中已有2名玩家使用与你相同的序列号.7   There are no more free slots in that game for your side6   你方在那场比赛中没有更多的免费槽位了E   This map has a %d player max.  The max includes human and AI players.A   这张地图有%d玩家上限. 上限包括人类和电脑玩家.   This may give the host   这可能会交给主机*   This product requires a 16bit pixel depth!!   此产品需要16位像素深度!   Tiberian Sun   泰伯利亚之日   Tiberian Sun BattleClans   泰伯利亚之日BattleClans   Tiberian Sun Disk %d   泰伯利亚之日光盘 %d   Tiberian Sun Players   泰伯利亚之日玩家   Tiberian Sun game channels   泰伯利亚之日游戏频道3   Tiberian Sun is unable to detect your CD ROM drive.7   泰伯利亚之日无法检测到您的CD ROM驱动器.�   Tiberian Sun requires %s version %d.%d or newer.

Please consult the read me for instructions on how to
obtain a newer version of %s.j   泰伯利亚之日需要 %s 版本%d.%d或更新.

请参考readme的了解如何获取
较新版本的%s./   Tiberian Sun will now restart to update itself.=   泰伯利亚之日现在将重新启动以进行自我更新.   Tiberium Lifeforms   泰伯生命体   Time allowed: %02d seconds   允许时间:%02d秒   Time of Day Transitions   一天中的时间转换   Time:%02d:%02d   时间:%02d:%02d   Time:%02d:%02d:%02d   时间:%02d:%02d:%02d   Tiny Map	   小地图   To %s:   致 %s:   To All:   致所有人:�   To start a BattleClan tournament game there needs to be an even number of people from two clans.  Everyone in the game must be in a clan.~   要开始BattleClan锦标赛游戏, 需要来自两个氏族的偶数玩家. 游戏中的每个人都必须属于一个氏族..   Toggle alliance with owner of selected object..   与选定对象的所有者切换联盟状态.*   Toggle follow state of selected object(s)."   切换选定对象的跟随状态.   Toggle power mode on / off.   打开/关闭电源模式.#   Toggle radar display mode on / off.!   切换雷达显示模式 开/关.   Toggle repair mode on / off.   打开/关闭修复模式.   Toggle sell mode on / off.   打开/关闭出售模式.(   Toggle waypoint placement mode on / off.#   打开/关闭路径点放置模式.   Tournament Game   锦标赛游戏   Tournament:
   锦标赛:  Tratos is being held in a hospital prison facility within this sector.  Avoid detection and rescue Tratos from the facility.  Once he is out, a transport will be sent in to evacuate him.  Once Tratos is clear, destroy all Nod forces in the area to prevent further experimentation.�   特拉托斯被藏在本区的一所监狱设施中, 潜入并救出他. 他出来之后, 我们会派一辆运输车来带他撤离. 特拉托斯安全之后, 摧毁该地区所有Nod部队以阻止他们继续实验.   Tundra   冻土   Two Player Only   仅限两名玩家-   Unable to find modem. Check power and cables.0   找不到调制解调器. 检查电源和电缆.A   Unable to join original Tiberian Sun game with Firestorm enabled.O   无法在火焰风暴开启的情况下加入原版泰伯利亚之日的游戏.+   Unable to play Direct Sound primary buffer.%   无法播放Direct Sound主缓冲区.#   Unable to play; scenario not found.   无法继续; 未找到场景.   Unable to read scenario!   无法加载场景!   Unit List Down   单位列表向下   Unit List PageDown   单位列表向下翻页   Unit List PageUp   单位列表向上翻页   Unit List Up   单位列表向上   Units   单位   Unknown Ping   未知的 Ping   Unknown Status   未知状态   Unlimited Game Length   无限游戏长度   Unranked	   未排名%   Unrecognized Direct Draw result code.&   无法识别的DirectDraw结果代码.   Unrevealed Terrain   未探索之地形�   Use the cyborg commando and his team to locate the bio-toxin tanker trucks.  Both trucks must reach the convoy point here if they are to arrive in time to aid you in your assault against the research facility.  GDI patrols are known to be in the area.�   使用生化尖兵来定位生物毒素油罐车. 两辆卡车必须到达护送点才能一起出发, 并引导你攻击研究设施. 情报显示, 在该地区附近还有GDI的巡逻队.*   User %s was kicked out of channel %s by %s   用户 %s 被 %s 踢出频道%s   User chat channels   用户聊天频道   User has find disabled   用户已禁用查找   User has pages disabled   用户已禁用页面   User is in channel %s   用户位于频道 %s 中   User isn't in any channels   用户不在任何频道中   User isn't logged in   用户未登录   User signed off!   用户已签名:   V.Large	   非常大0  Vega's base is secreted on an island in this sector.  Reaching it will be difficult, as there is only one overland access.  Your best chance of success lies in the use of amphibious APCs to land on the island and penetrate Vega's defenses.  Once on the island, destroy Vega's facility and command center.�   维加的基地在这里一个岛上. 要从陆上到达那里会很困难, 因为只有一条通道. 而你最好选择使用运兵车登陆岛屿并穿过维加的防御. 上岛之后, 立即摧毁维加的设施和指挥中心.	   Veinholes	   脉络孔   Very Abundant   非常丰富   Very Abundant Tiberium   非常丰富的泰矿   Very Abundant Water   非常丰富的水   Very Few	   非常少   Very Few Cities   非常少的城市   Very Few Cliffs   非常少的悬崖   Very Few Hills   非常少的山丘   Very Few Tiberium Fields   非常少的泰矿
   Very Heavy   非常厚重   Very Heavy Vegetation   非常厚重的植被	   Very High	   非常高   Very High Accessibility   非常高的可访问性   Very Low	   非常低   Very Low Accessibility   非常低的可访问性	   Very Many	   非常多   Very Scarce   非常稀缺   Very Scarce Tiberium   非常稀缺的泰矿   Very Scarce Water   非常稀缺的水   Very Sparse   非常稀疏   Very Sparse Vegetation   非常稀疏的植被   Video   显示   View Bookmark 1   查看书签 1   View Bookmark 2   查看书签 2   View Bookmark 3   查看书签 3   View Bookmark 4   查看书签 4   View bookmarked map position 1.   查看书签地图位置 1.   View bookmarked map position 2.   查看书签地图位置 2.   View bookmarked map position 3.   查看书签地图位置 3.   View bookmarked map position 4.   查看书签地图位置 4.   Voice   声音   WDT GDI Players   WDT GDI 玩家   WDT Nod Players   WDT Nod 玩家   Waiting for Call...   等待电话...(   Waiting for GO response - Please Wait...#   正在等待GO响应 - 请稍候...   Waiting for Opponent   等待对手-   Waiting for all players to enter the game....!   等待所有玩家进入游戏...   Waiting to Connect...   正在等待连接.../   Warning - Unable to create Direct Sound Object.(   警告 - 无法创建Direct Sound对象.7   Warning - Unable to create Direct Sound primary buffer..   警告 - 无法创建Direct Sound主缓冲区.7   Warning - Unable to set Direct Sound cooperative level..   警告 - 无法设置Direct Sound合作级别.I   Warning - Your sound card does not meet the product's audio requirements.4   警告 - 您的声卡不符合产品的音频要求.E   Warning - you are critically low on free disk space for saving games.7   警告 - 你的可用磁盘空间不足以保存游戏.n   Warning - you are critically low on free disk space for saving games. Do you want to play Tiberian Sun anyway?f   警告 - 用于保存游戏的可用磁盘空间严重不足. 你仍想继续玩泰伯利亚之日吗?   Warning: Ion Storm approaching.!   警告: 离子风暴即将来临.   Warning: Ion Storm here!   警告: 离子风暴来了!   Waypoint Mode   路径点模式  We have become aware of an imprisoned commander in this region who WAS loyal to Hassan.  Free him and his forces and they should be sympathetic to our cause -- and help in the capture of Hassan.  The commander may have information vital to my.......your movement.�   我们得知在这个地区有一个被囚禁的指挥官, 他曾忠于哈桑. 释放他和他的军队并加以利用, 这应该能帮助我们抓住哈桑. 这位指挥官可能有对我...你的事业至关重要.K  We must destroy GDI's new weapon.  They will, of course, build more in the future but it will buy us valuable time.  We know GDI is testing the Mammoth somewhere in this sector.  Use a chameleon spy to infiltrate a GDI comm center and locate the test site.  Your fighter prototype should be all you need to obliterate the nuisance.4  我们必须摧毁GDI的新武器. 虽然他们将来还会建造更多, 但这将为我们争取宝贵的时间. 我们知道GDI正在这个领域的某个地方测试猛犸机甲. 使用变色龙间谍渗透GDI通信中心并定位测试地点. 你的原型战斗机就是你消除麻烦所需要的一切.3  We suggest that the brotherhood should not suffer the indignations of the past.  In order to prevent history from repeating itself, you must steal the firing codes for GDI's ion cannon.    Paranoid security measures prevent GDI from storing the entire code in one place.  Therefore, use a chameleon spy to infiltrate three different comm centers.  Once we have the codes and the spy is safely evacuated, we will be able to use GDI's ion cannon against them in the final assault.  Unfortunately GDI will have to use the ion cannon once before we can use the codes.�  我们建议兄弟会不要再忍受过去的屈辱了. 为了防止历史重演, 你必须窃取GDI离子炮的发射代码. 以GDI的安全意识, 他们不会将代码存储在一个地方. 因此, 使用变色龙间谍渗透到三个不同的通信中心. 找到代码后立刻撤离间谍, 我们就可以在最后的攻击中使用GDI的离子炮来对付他们. 不幸的是, 必须先让GDI发射一次离子炮我们才能够使用代码.   Web Page   网页=   Would you like to launch your web browser to visit this page?+   您想启动web浏览器访问此页面吗?&   Would you like to replay this mission?   您想重玩此任务吗?   Yellow   黄色   Yes   是   You Are Victorious!   你胜利了!$   You are not in a Tiberian Sun squad.%   你不属于泰伯利亚之日小队.T   You can't make a channel with this name.  Try removing spaces and other punctuation.N   你不能用这个名字创建频道. 试着去掉空格和其他标点符号.W   You can't make a channel with this password. Try removing spaces and other punctuation.N   您无法使用此密码创建频道. 尝试删除空格和其他标点符号.D   You can't propose removing yourself. Click cancel to leave the game.8   你不能提议自己离开. 单击"取消"退出游戏.   You can't reject yourself!   你不能拒绝自己!5   You can't send a message when you're not in a channel,   当您不在频道中时, 无法发送消息<   You cannot change alliances in a World Domination Tour game.4   你不能在世界统治之旅游戏中改变结盟.   You cannot create this channel.   您无法创建此频道.0   You cannot kick a player from a tournament game.%   你不能在锦标赛中踢出玩家.8   You don't have a web browser associated with HTML files./   您没有与HTML文件相关联的web浏览器.g   You have not set your location. Click OK to continue anyway or cancel to go back and set your location.Z   您尚未设置地区. 单击"确定"继续, 或单击"取消"返回并设置您的地区.   You joined channel %s   你已加入频道 %s   You left channel %s   您离开了频道 %s*   You must be a channel operator to do this.1   您必须是频道运营商才能执行此操作..   You must be in a BattleClan to join this game.2   你必须在BattleClan中才能加入这个游戏.   You must enter a description!   您必须输入描述!   You must enter a name!   你必须输入一个名称!G   You must have an equal number of GDI and Nod players to start the game.@   你必须拥有相同数量的GDI和Nod玩家才能开始游戏.e  You must reach the medical colony in the region without being prematurely detected by GDI and forcing a base evacuation.  To prevent this, consider first destroying the 3 sensor towers protecting the base.  Our new artillery unit should be sufficient for the job, even in your hands.  Once inside the base, the capture of the mutant female should be simple.   你必须在不被GDI过早发现并迫使基地撤离的情况下到达该地区的医疗基地. 为了防止这种情况, 首先考虑破坏保护基座的3个传感器. 我们的新炮兵部队应该足以胜任这项工作. 一旦进入基地, 捕获那个女变种人应该很简单.   You must select a game!   你必须选择一个游戏!#   You must select a player to reject."   您必须选择要拒绝的玩家./   You must select a user to kick/ignore/ban them.6   你必须选择一个用户来踢/忽略/禁止他们.&   You need %d players to start the game.)   你还需要 %d 个玩家来开始游戏.*   You need to enter the same password twice.%   您需要输入相同的密码两次.'   You were kicked out of channel %s by %s   您被 %s 踢出了频道 %s0   You've been banned from Westwood Online until %s0   您已被禁止在 %s 之前访问Westwood网络$   You've been banned from this channel   您已被禁止进入此频道(   You've been disconnected from the server   您已与服务器断开连接`   You've been temporarily banned. Would you like to open your web browser to get more information?H   你被暂时封禁了. 您想打开web浏览器以获取更多信息吗?i   Your Serial number is currently in use.  Would you like to open your web browser to get more information?W   您的序列号当前正在使用中. 您想打开web浏览器以获取更多信息吗?�   Your account has been temporarily disabled.  Make sure the Email address you registered with is correct.  Would you like to open your web browser to get more information?�   您的帐户已被暂时禁用. 请确保您注册的电子邮件地址是正确的. 您想打开浏览器获取更多信息吗?   Your game name must be unique.%   您的游戏名称必须是唯一的.   Your game version is outdated.   您的游戏版本已经过时.   Your name must be unique.   你的名字必须是唯一的.-   Your password must be exactly 8 letters long.)   您的密码必须正好是8个字母长./   Your player name is blank, please enter a name.0   您的玩家名称为空, 请输入一个名称.�   Your serial number is associated with a product other than Tiberian Sun.  You must reinstall the game, specifying a valid Tiberian Sun serial number, to play online.�   您的序列号与泰伯利亚之日以外的产品相关联. 您必须重新安装游戏, 指定有效的泰伯利亚之日序列号, 才能游玩在线游戏.�   Your serial number was not found.  This is most likely due to a mistyped serial number during installation.  You must reinstall the game, specifying a valid serial number, to play online.�   找不到您的序列号. 这很可能是由于在安装过程中输入了错误的序列号. 您必须重新安装游戏并指定有效的序列号才能游玩在线游戏.   [%s's Game]   [%s 的游戏]   [EMPTY SLOT]   [空槽位]   [NONAME]   [无名氏]
   [OBSOLETE]   [过时]   a modified map.   修改后的地图.   an unfair advantage.   不公平的优势.   disconnected from the network.   与网络断开连接.1   disconnected from your internet service provider..   与您的互联网服务提供商断开连接.1   players don't elect to remove you from the game..+   玩家不会选择将你从游戏中移除.P   you can re-dial your provider and continue the game as normal provided the other    
ts_mission    K      A New Beginning   NOD 12A: 一个新的开始�  Another possible location of the Prototype Manufacturing Facility. Use the mutants to locate the position of the production facility. They must remain undetected. If Nod suspects enemy forces, they will cloak their production facility and deploy troops to destroy them. If the mutants can hide from the Nod troops for a short period, then Nod will assume the area is clear and uncloak the base. Once we record the location of the base, GDI Dropships will arrive with reinforcements.@@Objective One: Using Mutants you must locate the Prototype Manufacturing Facility.@@Objective Two: Once the facility is located reinforcements will be sent into help construct a base. You are to destroy the manufacturing facility at this time.�  原型制造设施的另一个可能位置. 利用变种人定位生产设施的位置. 变种人必须保持隐蔽. 如果Nod怀疑敌军存在, 他们将隐形设施并增加部队. 如果变种人能在短时间内躲避Nod部队, Nod将认为区域安全并解除设施隐形. 记录设施位置后, GDI空降兵将携援军抵达.@@目标一: 利用变种人定位原型制造设施.@@目标二: 一旦找到设施, 建立基地并摧毁设施.o  BE ADVISED: Kane is determined to destroy you. He knows the Kodiak cannot lift off during an ion storm and has chosen this moment to attack. The Kodiak must be protected until the storm abates. The storm will interfere with certain types of equipment so expect some malfunction.@@Objective One: Protect the Kodiak at all costs.@@Objective Two: Destroy all Nod forces.+  注意: 凯恩决心消灭你. 他知道离子风暴期间科迪亚克无法起飞, 于是选择此时发动攻击. 你必须保护科迪亚克直到风暴结束. 风暴会干扰某些设备, 预计会出现故障.@@目标一: 不惜一切代价保护科迪亚克.@@目标二: 消灭所有Nod部队.   Blackout   NOD 04B: 灯火管制   Capture Hammerfest Base#   GDI 07: 夺回哈默菲斯特基地   Capture Jake McNeil"   NOD 11: 抓获杰克·麦克尼尔   Capture Train Station   GDI 03B: 占领火车站   Capture Umagon   NOD 06A: 逮捕乌玛贡�  Control of the mutants is in our grasp. Their headquarters is located to the north of your drop-off position. The units you will need to implicate GDI in this deception can be obtained by capturing the rest of the GDI base that you will start in. Do not mar the Brotherhoods name any further. Allow the blame to fall squarely upon Solomon's shoulders.@@Objective One: Capture the enemy Construction Yard awaiting you.@@Objective Two: Use GDI units to destroy the mutant's base.  我们将掌握变种人的控制权. 他们的总部在你的北边, 你需要通过占领GDI基地获得兵力补给. 不要再玷污兄弟会的名声, 让责任全部落到所罗门头上. @@目标一: 占领敌方建造厂.@@目标二: 使用GDI部队摧毁变种人基地.   Defend Crash Site   GDI 04: 防守坠毁现场   Destroy Chemical Missile Plant!   GDI 09A: 摧毁化学导弹工厂   Destroy Chemical Supply   GDI 09B: 切断化学品供应   Destroy GDI Research Facility   NOD 07A: 摧毁GDI研究设施   Destroy Mammoth Mk.II Prototype#   NOD 10: 摧毁猛犸机甲原型机   Destroy Prototype Facility    GDI 10: 摧毁原型制造设施   Destroy Radar Array   GDI 05B: 摧毁雷达阵列   Destroy Vega's Base   GDI 06A: 摧毁维加的基地   Destroy Vega's Dam   GDI 06B: 摧毁维加的水坝�   Destroy the three relay stations and the radar array to blackout Nod's sensor net. This will make rescuing Tratos easier, as Nod will not be as quick to detect you.@@Objective One: Destroy the three relay stations.@@Objective Two: Destroy the radar array.�   摧毁三座中继站和雷达阵列以瘫痪Nod的传感网络. 这将使营救特拉托斯变得更加容易, 因为Nod将无法迅速发现你.@@目标一: 摧毁三座中继站. @@目标二: 摧毁雷达阵列.   Detroy Hassan's Temple   NOD 03A: 摧毁哈桑的神殿�  Emergency transmissions from GDI forces in this region indicate that Phoenix Base is under attack from Nod troops. It is imperative that the base be restored by building a Tiberium Refinery and a Barracks. Once the base is functional, all Nod forces in the area must be destroyed.@@Objective One: Build a Tiberium Refinery.@@Objective Two: Build a Barracks.@@Objective Three: Destroy all Nod forces.b  来自该区域GDI部队的紧急通讯显示, 费城基地正遭到Nod部队的攻击. 当务之急是通过建造一座泰矿精炼厂和一个兵营来恢复基地运作. 一旦基地恢复正常, 你必须消灭该区域内的所有Nod部队.@@目标一: 建造一座泰矿精炼厂.@@目标二: 建造一个兵营.@@目标三: 消灭所有Nod部队.   Escort Bio-toxin Trucks!   NOD 07B: 护送生物毒素卡车   Establish Nod Presence   建立Nod驻防队   Eviction Notice   NOD 04A: 驱逐通知   Final Conflict   GDI 12: 最终冲突   Free Rebel Commander   NOD 03B: 释放叛军指挥官�  GDI forces in this sector have found something unusual and large that crashed nearby. Nod has taken an intense interest in whatever it is, so naturally we are interested as well. Locate the object from the reports and capture any Nod Technology Centers in the area that might have uncovered clues as to the identity of the object.@@Objective One: Locate the Crash Site.@@Objective Two: Capture any Nod Technology Centers.  该区域的GDI部队发现了一个奇怪的坠落物. Nod对此表现出极大兴趣, 因此我们也自然不能忽视. 你需要找到该坠落物, 并占领区域内可能揭示其身份线索的Nod科技中心.@@目标一: 找到坠毁地点.@@目标二: 占领Nod科技中心.[  GDI has secured the Holy Ground the temple rests on. Your objective is simple, locate it and remove the GDI incursion. They are not expecting any Nod forces, so the element of surprise is yours. The temple and its knowledge must remain intact. One vision, One purpose!@@Object One: Locate the Temple of Nod.@@Objective Two: Destroy all GDI forces.1  GDI已经占领了神殿所在的圣地. 你的任务很简单, 找到它并消灭GDI入侵者. 他们未预料到会有Nod部队出现, 因此你拥有出其不意的优势. 神殿及其知识必须保持完整. @唯有信念, 唯有使命!@@目标一: 找到Nod神殿.@@目标二: 消灭所有GDI部队.�  GDI has stored the firing codes for its Ion Cannon in three separate Comm centers. The centers are isolated in a valley and poorly guarded. We do not have the forces available for a full-scale assault. However, a small infiltration team led by the Chameleon Spy has a reasonable chance of success. Once the Spy has the codes, he must be evacuated safely.@@Objective One: Infiltrate the Comm centers and steal the codes.@@Objective Two: Evacuate the Chameleon Spy.y  GDI将离子炮的发射代码分别存放在三座通讯中心中. 这些中心被隔离在一个山谷中, 戒备森严. 我们没有足够兵力发动全面进攻. 然而, 由变色龙间谍率领的小型渗透小队有成功的机会. 一旦间谍获取代码, 必须确保他安全撤离.@@目标一: 潜入通讯中心并窃取代码. @@目标二: 撤离变色龙间谍.  GDI is set to test the prototype of their new weapon, the Mammoth Mark II. It is vital that we sabotage their production of this monster as soon as possible. Before we can do that however, we need to know where the test is being held. Send a Chameleon Spy into one of the Radar Facilities. The coordinates to the testing ground should be stored there. Be careful of the patrols in the area - we have only one spy available. Once we have the location of the test, construct a base and destroy the prototype. You now have access to the new Banshee aircraft, which should prove useful. Destroying the remainder of the GDI base is at your discretion, but the Mammoth MUST be destroyed.@@Objective One: Spy on one of the GDI Comm Centers.@@Objective Two: Destroy the Mammoth Mark II prototype.�  GDI准备测试他们的新型武器原型 - 猛犸二型机甲. 这头怪物的生产必须尽快被破坏. 然而在那之前, 我们需要知道测试地点的位置. 派出一名变色龙间谍潜入一座雷达设施. 测试场的坐标应该存储在那里. 要小心该区域的巡逻队 - 我们只有一名间谍可用. 一旦获得测试地点, 立即建立基地并摧毁该原型机. 你现在已获得新型单位"女妖"战机的使用权限, 它应当会非常有用. 是否摧毁GDI基地的其余部分由你决定, 但猛犸必须被摧毁.@@目标一: 潜入一座GDI通讯中心进行侦查. @@目标二: 摧毁猛犸二型原型机.�  Hammerfest base has been overrun by Nod troops. The Firestorm walls block direct approach, so another route must be found back into the complex. Using hover MLRS and waterways for access, find a way back to the GDI base and re-capture it. Once the base is back in GDI hands, destroy all Nod forces in the area.@@Objective One: Find a way back to the GDI base.@@Objective Two: Re-capture the base with engineers.@@Objective Three: Destroy all Nod forces in the area.�  哈默菲斯特基地已被Nod部队攻占. 火焰风暴墙阻挡了正面通路, 必须另寻路径进入基地. 利用悬浮多管火箭发射车从水路进入, 设法返回GDI基地并重新夺回控制权. 一旦基地重归GDI之手, 消灭该区域内的所有Nod部队.@@目标一: 寻找返回GDI基地的路径.@@目标二: 用工程师重新夺回基地.@@目标三: 消灭该区域内的所有Nod部队.=  Hassan is determined to stop you at any cost. He has pursued us back to a small base near his HQ. We must fend off his assault and build a Tiberium Refinery so we have the means to strike back.@@Objective One: Get production online by building a Tiberium Refinery.@@Objective Two: Destroy all of Hassan's Elite Guard..  哈桑决心不惜一切代价阻止你. 他已经追击我们至其总部附近的一个小型基地. 我们必须抵挡住他的进攻, 并建造一座泰矿精炼厂, 以便具备反击的能力.@@目标一: 建造一座泰矿精炼厂以恢复生产. @@目标二: 消灭哈桑的所有精锐卫队.�  Hassan spreads his propaganda to the Brotherhood through a nearby TV station. With the Brotherhood in chaos, the opportunity to divide Hassan from his followers presents itself. Capture the TV station and those once loyal to Kane's technology of peace will return to the fold. And as for Hassan's pathetic guards - crush them.@@Objective One: Capture the TV station to the east.@@Objective Two: Destroy Hassan's Elite Guard.d  哈桑正在通过附近的电视台向兄弟会传播他的思想. 如今兄弟会陷入混乱, 正是分裂哈桑与其追随者的好时机. 占领这座电视台, 那些曾忠于凯恩"和平科技"的人将重归麾下. 至于哈桑的那些可怜的卫兵 - 粉碎他们.@@目标一: 占领东边的电视台.@@目标二: 消灭哈桑的精锐卫队.�  If the upcoming GDI attack on the missile sites is to succeed, C4 must be planted at all six power stations. The power grid is well protected, but the train should carry the demolition team and the mutants through the gates and past the guards. If Nod forces discover the demolition team and sound the alert, take out the power plants by any means available.@@Objective One: Plant C4 at the power plants.>  为了GDI对导弹基地的进攻取得成功, 必须在全部六座发电站安装C4炸药. 电力网络防守严密, 不过火车应该能将爆破小组和变种人送入大门. 如果Nod部队发现了爆破小组并发出警报, 就无论一切手段摧毁这些发电站. @@目标一: 在发电站安放C4炸药.   Illegal Data Transfer   NOD 12B: 非法数据传输�  Impulses scanned from signatures emanating from Cairo suggest Kane will launch his world-altering missile within hours. You must destroy the Pyramid Temple before he has a chance to launch. There are no other strategies.@@Objective One: Clear the zone for MCV Dropship deployment.@@Objective Two: Destroy the ICBM launchers.@@Objective Three: Destroy the Pyramid Temple.@@Objective Four: Destroy all Nod forces.G  从开罗发出的信号表明, 凯恩将在几小时内发射他那足以改变世界的导弹. 你必须在他发射之前摧毁金字塔神殿. 没有其他的策略.@@目标一: 为MCV的部署清理区域.@@目标二: 摧毁洲际弹道导弹发射器.@@目标三: 摧毁金字塔神殿.@@目标四: 摧毁所有Nod部队.�  In order for our ICBMs to shoot down the Philadelphia, they must be able to triangulate the station's position. Our spies have placed beacons at the optimal deployment locations. Once the launchers have been moved to the beacons, the station's fate is sealed and the Temple of Nod may be built. Move with all due haste. If the Philadelphia is able to complete three orbits, it will lock onto our position and destroy Kane's plans.@@Objective One: Deploy ICBM launchers at the three beacons.�  为了让我们的洲际弹道导弹击落费城空间站, 必须能够三角定位该空间站的位置. 我们的间谍已在最佳位置放置了信标. 一旦我们的发射器在信标处就位, 空间站的命运就注定了, Nod神殿也将会建成. 务必迅速行动, 如果空间站锁定了我方位置, 凯恩的计划将会遭到致命打击.@@目标一: 在三个信标处部署洲际弹道导弹发射器.?  It is imperative that you prevent the train carrying the crystals from reaching the Nod base. Recent ice melts in the region have washed out the only train bridge. However, Nod engineers are on their way to repair it, so you must move quickly. If you can get to the train before the bridge is repaired, we can recover the crystals with little trouble. Otherwise, we will have to assault the Nod base to reclaim the crystals. Remember, to stop the train, you must destroy the locomotive, not the cars, but the cargo car holds the crystals.@@Objective One: Locate the train and destroy the locomotive before Nod engineers repair the bridge. The cargo car holds the crystals.@@Objective Two: If the bridge is repaired and the train successfully reaches the Nod base, then you must locate and destroy this base to recover the crystals.X  你必须阻止运载水晶的火车到达Nod基地. 最近该地区的冰融化冲毁了唯一的火车桥. 然而, Nod的工程师正在修理它的路上, 所以你必须迅速行动. 如果你能在桥修好之前找到火车, 我们就能轻而易举地取回水晶. 否则, 我们就得攻击Nod基地夺回水晶. 记住, 要让火车停下来, 你必须摧毁火车头, 不是车厢, 特别是装有水晶的车厢.@@目标一: 在Nod工程师修理桥梁之前摧毁火车头.@@目标二: 如果桥被修复并且火车成功到达Nod基地, 那么你必须摧毁这个基地来夺回水晶.-  Jake McNeil, brother of one of GDI's commanders, will be leading an inspection tour to a small GDI outpost in this area. His knowledge of GDI activities could be of great benefit to Nod's cause. Capture the GDI outpost with engineers, then disguise the base as GDI's and wait for Jake to make his inspection. When the signal is given, use the Toxin soldiers provided to "persuade" Jake to join Nod's forces. Once he is under our influence, EVAC him at the designated site.@@@Be very careful not to alert GDI until we are ready to strike. If they detect Nod forces in the area, they will surely try to evacuate Jake. If GDI is alerted, be sure to get to Jake before he can leave the area.@@Objective One: Capture the GDI outpost.@@Objective Two: Capture Jake.@@Objective Three: EVAC Jake at the specified location.�  杰克·麦克尼尔是GDI一名指挥官的兄弟, 他将带领一支巡查队伍前往GDI在这个地区的一个小前哨. 他对GDI的了解对Nod的事业大有裨益. 用工程师占领GDI的前哨, 然后把基地伪装成GDI的基地, 等待杰克到来. 当信号发出时, 使用毒素步兵来"说服"杰克加入Nod部队. 一旦他被我们"说服", 就把他撤离到指定地点.@@@在我们准备好之前, 要小心不要惊扰GDI. 如果他们发现这是陷阱, 肯定会设法撤离杰克, 如果变成这样, 一定要在杰克逃跑之前抓住他.@@目标一: 占领GDI前哨.@@目标二: 抓住杰克·麦克尼尔.@@目标三: 在指定地点撤离杰克.   Mine Power Grid   GDI 09C: 摧毁矿场电网�  Nod forces were recently forced out of this area. However, spies report that the Nod bio-toxin facility has not yet been destroyed by GDI troops. The Cyborg Commando and his team should be able to slip through the main GDI force and recover two tankers full of bio-toxin - provided we act quickly.@@Objective One: Locate the bio-toxin trucks.@@Objective Two: Escort the trucks to the checkpoint east of the base.B  Nod部队最近被迫撤出这个地区. 然而, 间谍报告称, Nod生物毒素设施尚未被GDI部队摧毁. 只要我们迅速采取行动, 生化尖兵应该能够穿过GDI部队, 回收两辆装满生物毒素的卡车.@@目标一: 定位生物毒素运输车.@@目标二:护送卡车前往基地以东的检查站.%  Nod has positioned a supply base in the area near a civilian train station. We can use the train and supplies to infiltrate the larger Nod base to the east. Avoiding patrols where possible and destroy all the Nod structures in the area. Once the area is secure, capture the train station for our use. DO NOT destroy the station or the train, as they are vital to our plans. Engineers and other reinforcements are available, but not unlimited - do not waste them.@@Objective One: Destroy all Nod structures.@@Objective Two: Capture the train station.�  Nod在民用火车站附近的地区建立了一个补给基地. 我们可以利用火车渗透到东部更大的Nod基地. 尽可能避免与巡逻队接触, 并摧毁该地区的所有Nod建筑. 一旦该地区安全, 占领火车站供我们使用. 不要破坏车站或火车,  因为它们对我们的计划至关重要. 工程师和其他增援部队是可用的, 但不是无限的 - 不要浪费.@@目标一: 摧毁所有Nod建筑.@@目标二: 占领火车站.�  Nod is experimenting on mutant survivors at a facility in this sector. Among them is Tratos, leader of the mutants. Using Umagon's strike team, rescue Tratos from imprisonment and EVAC him at the specified site. Once complete, move in with GDI forces and destroy the Nod base and the prison test facility.@@Objective One: Rescue Tratos from prison.@@Objective Two: EVAC Tratos at specified site.@@Objective Three: Destroy the Nod base and test facility.�  Nod正在该地区的一个设施对变种人存者进行实验. 其中包括变种人的领袖特拉托斯. 使用乌玛贡的突击队, 将特拉托斯从医院中救出, 并在指定地点将其撤离. 完成后, 与GDI部队一起行动, 摧毁Nod基地和相关设施.@@目标一: 从医院中营救特拉托斯.@@目标二: 在指定地点撤离特拉托斯.@@目标三: 摧毁Nod基地和相关设施.|  Nod's main chemical missile plant is located in this area. It is responsible for the large amount of Tiberium poisoning and accelerated mutations of wildlife in the surrounding areas. Destroying this facility will prevent Nod from furthering the acceleration of Tiberium poisoning on the planet.@@Objective One: Destroy Nod's missile silos.@@Objective Two: Destroy all Nod forces.#  Nod的主要化学导弹工厂就在这个地区. 该工厂是周边地区大量泰伯利亚污染和野生动植物加速变异的根源. 摧毁这个设施将阻止Nod进一步加剧泰伯利亚对地球的污染.@@目标一: 摧毁Nod的导弹发射井.@@目标二: 摧毁所有Nod部队.�  One of two possible locations of the Prototype Manufacturing Facility. Use the mutants to locate the position of the production facility. The mutants must remain undetected. If Nod suspects enemy forces in the area, they will cloak the facility and deploy troops to destroy them. If the mutants can hide from the Nod troops for a short period, the base will assume the area is clear and uncloak. Once we record the location of the base, GDI Dropships will arrive with reinforcements.@@Objective One: Using mutants you must locate the Prototype Manufacturing Facility.@@Objective Two: Once the facility is located, reinforcements will be sent in to help construct a base. You are to destroy the Manufacturing Facility at this time.�  原型制造工厂的两个可能地点之一. 利用变种人定位工厂的位置. 变种人必须不被发现. 如果Nod怀疑该地区有敌军, 他们会隐形设施并派兵摧毁敌人. 如果变种人能躲过Nod的部队一段时间, 基地就会认为这片区域已安全并解除隐形. 一旦我们得到基地的位置, GDI的援军就会到达. @@目标一: 利用变种人定位原型制造设施.@@目标二: 摧毁原型制造工厂.   Protect Waste Convoys#   NOD 09: 保护泰矿物质运输车   Reestablish Nod Presence   NOD 09: 恢复NOD驻扎   Reinforce Phoenix Base   GDI 01: 增援费城基地   Rescue Prisoners!   GDI 09D: 营救被遗忘者囚犯   Rescue Tratos   GDI 05A: 营救特拉托斯   Retaliation   NOD 02: 报复   Retrieve Disrupter Crystals   GDI 08: 夺回声波晶体   Salvage Operation   NOD 05: 打捞作业   Secure Crash Site   GDI 03A: 清空坠毁现场   Secure The Region   GDI 02: 确保区域安全   Sheep's Clothing   NOD 06B: 披着羊皮的狼K  Taking out this weak position of GDI forces will allow us to reclaim our Sarajevo temple without interruption. Move in under the cover of an ion storm - while GDI's communications will be down. Take out the Radar Facility before the storm abates.@@Objective One: Locate and destroy the GDI Radar Facility before the ion storm ends.�   摧毁GDI这一薄弱据点, 将使我们能够顺利收复萨拉热窝神殿. 利用离子风暴作为掩护行动 - 此时GDI的通讯将中断. 在风暴结束前摧毁雷达设施.@@目标一: 在离子风暴结束前找到并摧毁GDI雷达设施.�  The Cyborg Commando has been sent in to retrieve you. Once free, rendezvous with your rescue team to the south. Use them to locate and free Oxanna. She will soon be transported to the main GDI facility, optimal chances for success rely on obtaining her before she is transported. After she has been freed, commandeer a GDI transport to make your escape.@@Objective One: Locate and free Oxanna.@@Objective Two: Steal a GDI transport to make an escape.@  生化尖兵前去营救你. 获救后, 与救援队会合. 利用他们寻找并救出奥克斯安娜. 她很快将被送往GDI主基地, 成功的关键是要在她被转移前救出她. 救出后, 夺取一辆GDI运输机逃离. @@目标一: 找到并救出奥克斯安娜.@@目标二: 夺取GDI运输机进行撤离.K  The Infidel, Hassan, has been tracked to this region of Cairo. Build a base and eliminate this would-be pharaoh, the pretender to Kane's throne.@@Objective One: Cross the bridge and destroy the enemies on the far side.@@Objective Two: Deploy your MCV and begin building a base.@@Objective Three: Locate and destroy Hassan's Temple.  异教徒哈桑已被追踪到开罗的这一地区. 建立基地, 消灭这个妄图篡夺凯恩王位的冒牌货.@@目标一: 穿过桥梁, 消灭桥对岸的敌人.@@目标二: 部署你的基地车并开始建设基地.@@目标三: 找到并摧毁哈桑的神殿.   The Messiah Returns   NOD 01: 弥赛亚归来�  The Nod base in this sector has been overrun by Tiberium life forms. Weedeaters have proven to be effective against the Tiberium creatures, but we must move reinforcements in quickly before the base is completely destroyed. Once the situation has been stabilized, the GDI base in the area must be eliminated.@@Objective One: Locate and secure the old base.@@Objective Two: Destroy the GDI base.  该地区的Nod基地已被泰伯生命体占领, 回收者对它们效果显著, 但我们必须在基地被完全摧毁之前迅速派遣增援部队. 局势稳定下来后, 必须消除该地区的GDI基地.@@目标一: 找到并保护旧基地.@@目标二: 摧毁GDI基地.g  The Nod forces that attacked Phoenix Base have been traced back to a small base in this sector. Orders received from GDI Command state that the Nod base must be destroyed. However, there is a significant civilian population in the immediate area that must be evacuated by ORCA Transport before the fighting gets too heavy. Before the Transports can safely land, all seven SAM sites must be destroyed. Once the civilians have been evacuated, the Nod base can be destroyed.@@Objective One: Deploy the M.C.V. and begin building a base.@@Objective Two: Destroy all Nod SAM sites.@@Objective Three: Destroy the Nod base.�  袭击费城基地的Nod部队已经追溯到这个区域的一个小基地. GDI指挥部下令必须摧毁该Nod基地. 但该区域内有大量平民, 必须在战斗加剧前由奥卡运输机撤离. 在运输机能够安全着陆之前, 必须摧毁七个萨姆飞弹发射阵地. 平民被疏散后, 就可以放心地摧毁Nod基地.@@目标一: 部署基地车开始建造基地.@@目标二: 摧毁所有萨姆飞弹发射台. @@目标三: 摧毁Nod基地.�  The alien craft is located in this region. FIND IT! The area is infested with GDI, so stealth would be to your advantage. Once the craft is located get an engineer inside to retrieve the Tacitus. And, should you encounter Vega's forces - consider them expendable.@@Objective One: Locate the crashed UFO and retrieve Kane's artifacts.@@Objective Two: Stop the transport of the Tacitus at all costs.p  外星飞船位于这个地区, 找到它! 这个地区到处都是GDI, 所以隐形对你十分有利. 一旦找到飞船, 让一名工程师进去取回塔西佗. 另外, 如果你遇到维加的部队, 放心用, 他们是可以牺牲的.@@目标一: 找到坠毁的不明飞行物并为凯恩取回塔西佗.@@目标二: 不惜一切代价阻止塔西佗的运输.'  The hydroelectric dams in this area provide Vega's island fortress with almost limitless power. Destroying the dams will seriously cripple Vega's perimeter defenses and allow GDI to bring more weapons to bear against Vega's base.@@The dams are heavily fortified, so attacking them directly is not the best option. Surveillance indicates the key to destroying the dams lies in the destruction of two regulator stations. Without them, the dams' generators will overload and the dams will self destruct.@@Objective One: Destroy the dams any way possible.�  该地区的水力发电大坝为维加岛的堡垒提供了几乎无限的电力. 摧毁水坝将严重削弱维加的周边防御, 使GDI能动用更多武器攻击维加基地.@@大坝防御严密, 因此直接攻击它们不是最好的选择. 侦察显示, 摧毁大坝的关键在于摧毁两个调节站. 没有它们, 大坝的发电机将会过载, 导致大坝自毁.@@目标一: 尽一切可能摧毁水坝.U  The mutant female may be trying to reach the underground railway system located in New Detroit. Move in and control the station before she arrives. If she boards the train then it must be stopped. This may be our last chance at capturing the abomination.@@Objective One: Locate the train station in the area and capture it before Umagon flies in and boards the train to escape into the underground.@Objective Two: If Umagon boards the train before you have captured the station then you must stop the train before it leaves the region. Destroy the locomotive and we will be able to capture Umagon.�  那名女性变种人可能正试图前往新底特律的地下铁路系统. 在她抵达之前, 赶往并控制车站. 如果她登上火车，必须将其拦下. 这也许是我们抓住这个异类的最后机会. @@目标一: 在乌玛贡登上火车之前, 找到该区域的火车站并将其占领. @@目标二: 如果在你占领车站之前乌玛贡已登上火车, 则必须在火车离开该地区前将其拦截并抓捕乌玛贡.�  The research facility in this sector must be destroyed before the GDI scientists perfect their Tiberium reduction technology. If Nod forces are to establish a base in the area, the GDI patrols must be eliminated. The mutants may prove to be useful allies.@@Objective One: Contact the mutants@@Objective Two: Clear GDI forces away from the tunnel and main road.@@Objective Three: Locate the research facility.@Objective Four: Destroy the research facility.j  在GDI科学家完善他们的泰伯利亚清除技术之前, 必须摧毁本区域的研究设施. 若Nod部队要在此地建立基地, 必须清除GDI的巡逻部队. 变种人或许能成为有用的盟友. @@目标一: 与变种人接触. @@目标二: 清除隧道和主干道上的GDI部队. @@目标三: 找到研究设施.@@目标四: 摧毁研究设施.�  The road through this sector is a vital supply link. If a foothold is firmly established and a Tiberium Waste Facility is built, Nod chemical missiles can be launched from the region. The GDI base in the area has no defense against the missiles, and can be destroyed at your leisure once the waste convoys start arriving.@@Objective One: Establish a base and build a Tiberium Waste Facility@@Objective Two: Destroy the GDI base.R  本区域是至关重要的补给通道. 如果能在此牢牢建立据点并建造一座泰矿物质回收厂, Nod就能从该地区发射化学导弹. 该区域的GDI基地对此毫无防御, 一旦运输车抵达, 你可以随时将GDI摧毁.@@目标一: 建立基地并建造一座泰矿物质回收厂. @@目标二：摧毁GDI基地./  This chemical supply station is providing vast quantities of Tiberium toxins to a number of Nod research programs in the area. Destroying this site will seriously hinder further Nod research, and prevent this base from transporting reinforcements to others in the sector.@@Intelligence reports advise caution when near any of the chemical tanks and facilities, as the toxins contained within are highly corrosive and equally deadly to soldiers and vehicles.@@Objective One: Find a suitable location for a base. Objective Two: Destroy the Nod Chemical station.�  该化学补给站正向本区域多个Nod研究项目提供大量泰伯利亚毒素. 摧毁此地将严重阻碍Nod的后续研究, 并阻止该基地向本区其他地点输送援军. @@情报提醒: 靠近任何化学罐体或设施时务必小心, 其中的毒素具有极强腐蚀性, 对士兵和载具都同样致命.@@目标一: 寻找合适地点建立基地.@@目标二: 摧毁Nod化学补给站.�  Umagon has requested help to rescue her people from a Nod prison. The prison is located on an island to the east. Nod has a strong force in the area, both in outposts and spread through the nearby city. We have limited resources and no reinforcements are available, so avoiding patrols is vital to your success. Umagon has a team in the area already - if you can find them, they may assist you. Make your way to the prison and release the hostages. Once the prison is secure, we will send a transport to evacuate Umagon's people. There may be SAM sites nearby, so make sure the way is clear for the transport.@@Objective One: Locate the Nod prison.@@Objective Two: Release and evacuate the prisoners.J  乌玛贡请求协助营救她的族人, 他们被关押在东边的一座Nod监狱中. Nod在该区域部署了大量兵力, 无论是在前哨还是在附近的市区, 我们的资源有限, 且没有增援部队, 因此需要尽可能避开巡逻队. 乌玛贡已有一支小队在该区域, 如果你能找到他们, 他们可能会提供帮助. 前往监狱并释放人质. 一旦监狱被控制, 我们将派遣运输机撤离乌玛贡的族人. 附近可能存在地对空导弹阵地, 请确保运输路径安全. @@目标一: 找到Nod监狱.@@目标二: 释放并撤离人质.�  Vega's base of operations is in the area. It is heavily guarded by SAM sites, and a secondary outpost provides reinforcements. Destroy all Nod forces in the area, but capture Vega's Pyramid intact - there is information there that we can use. You will have only limited troops until the SAM sites are neutralized one way or another.@@Objective One: Destroy the Nod base.@@Objective Two: Capture Vega's Pyramid.|  维加的作战基地位于此区域, 受到地对空导弹阵地的严密防护, 另有一个次级前哨提供增援. 消灭该区域内所有Nod部队, 但要完整地占领维加的金字塔 - 其中包含我们可利用的重要情报. 在地对空导弹阵地被清除之前, 你只能使用有限的部队.@@目标一: 摧毁Nod基地.@@目标二: 夺取维加的金字塔.   Villainess in Distress   NOD 08: 困境中的恶兽8  We have become aware of an imprisoned commander in this region who WAS loyal to Hassan. Free him and his forces and they should be sympathetic to our cause - and help in the capture of Hassan. The commander may have information vital to Hassan's movement.@@Objective One: Locate and free the Rebel Nod Commander.  我们得知该区域中关押着一名曾效忠于哈桑的指挥官. 释放他和他的部队, 他们应该会支持我们的事业, 并协助我们逮捕哈桑. 该指挥官可能掌握关于哈桑行动的重要情报.@@目标一: 找到并释放指挥官.   Weather the Storm   GDI 11: 挺过风暴  Whatever is contained in this craft, it is apparent that Nod doesn't want GDI to have it. Protect the crashed UFO until GDI reinforcements can arrive to fortify the area.@@Objective One: Survive until reinforcements can arrive.@@Objective Two: Prevent Nod from destroying the UFO.�   无论这艘飞船中装载着什么, 很明显Nod不希望GDI得到它. 在GDI援军抵达并加固该区域之前, 保护这艘坠毁的UFO.@@目标一: 坚持战线直到援军抵达.@@目标二: 阻止Nod摧毁UFO.E  You must reach the medical colony in the region without being prematurely detected by GDI and forcing a base evacuation. To prevent this, consider first destroying the three sensor towers protecting the base. Our new artillery unit should be sufficient for the job. Once inside the base, the capture of the mutant female should be easy.@@Objective One: Find and destroy the GDI sensor towers without getting too close and getting detected by them.@@Objective Two: Once the towers are destroyed, move on the base and capture the medical colony before Umagon, the Mutant, can escape.�  你必须在被GDI发现之前到达该地区的医疗殖民地. 为防止被提前发现, 建议优先摧毁保护基地的三座感应塔. 我们新的炮兵单位应该可以完成这项任务. 一旦进入基地, 要捕获那名女性变种人将变得轻而易举. @@目标一: 在不被发现的情况下, 找到并摧毁GDI的感应塔.@@目标二: 在变种人乌玛贡逃脱之前, 向基地推进到并占领医疗殖民地.ts_tutorial    �      ****BROADCASTING****   ****广播中****   Alert! GDI presence detected!   警报! 检测到GDI存在!    Alert! Prison break in progress!   警报! 囚犯们正在越狱!   BATTLEFIELD CONTROL ESTABLISHED   已建立战场控制!   Base perimeter has been breached!   基地外围已被攻破!2   Beware Tiberium is lethal to unprotected infantry..   小心泰矿对无保护的步兵是致命的.'   Build more infantry to defend the base!%   建造更多的步兵来保卫基地!   Bullet train departing.   火车出发了.�   CABAL: During the Ion Storm their Radar/Communications will be down. Now is the opportune time to hit them before the storm abates.|   CABAL: 在离子风暴期间, 他们的雷达/通讯将会中断. 现在是在风暴减弱之前袭击他们的最佳时机.]   CABAL: Establish a foothold on the far side of this bridge and an MCV will be sent in to you.L   CABAL: 在这座桥的另一边建立一个防线, 届时将派遣MCV支援.�   CABAL: Find and capture the train station before Umagon arrives. If she manages to make it onto a train then destroy it before she can escape.x   CABAL: 在乌玛贡到达之前找到并占领火车站. 如果她成功登上了火车那就在她逃脱之前摧毁它2   CABAL: GDI Communications have been reestablished.   GDI通讯已经重建.B   CABAL: General Vega, the generators are online.  SAM sites active.J   CABAL: 维加将军, 发生器已经启动. 萨姆飞弹发射台已激活M   CABAL: General Vega, the secondary generators will come online in 20 minutes.>   CABAL: 维加将军, 第二台发生器将在20分钟内启动:   CABAL: Hassan's Base has been alerted. Attack is imminent.9   CABAL: 哈桑基地已经收到警报, 攻击即将开始(   CABAL: MCV has arrived to the southeast."   CABAL: MCV已经到达东南方向.   CABAL: Philadelphia orbit tracking commencing!#   CABAL: 开始跟踪空间站轨道!#   CABAL: Slavik lost, mission failed.'   CABAL: 失去斯拉维克, 任务失败S   CABAL: With the train destroyed Umagon will be stranded.  Find her and capture her.2   CABAL: 火车已拦截, 乌玛贡被困, 抓住她   CAUTION: THIN ICE.   注意: 薄冰W   Captured Commander: All right! Now get me to your drop-off site and into the evac unit.E   被俘指挥官: 好吧! 现在带我去你的空投点, 送我撤离   Civilian city is under attack!   平民城市遭到攻击!.   Clear the zone for M.C.V. dropship deployment!   为MCV运输机清空区域!   Codes located.   代码已定位   Convoy destroyed.   已摧毁车队;   Current weapon range insufficient. Weapon drop in progress.,   当前武器射程不足. 正在投放武器7   Deploy the M.C.V. by double left clicking on the M.C.V.   通过双击左键来部署MCVH   Destroy the 7 SAM sites on the ridge to clear the way for our dropships.N   摧毁山脊上的7个萨姆飞弹发射台, 为我们的运输机扫清道路   Detonate C4 when ready.   准备好后引爆C4炸药   Down with Hassan!!!   打倒哈桑!!!+   ESTABLISHING BATTLEFIELD CONTROL - Standby!"   作战控制连接中 - 请稍后!j   EVA: Alert! The bridge has been fixed and the Nod train is moving to its final destination within the baseN   EVA: 警告! 桥梁已经修好, Nod列车正驶向基地内的最终目的地[   EVA: GDI reinforcements have arrived. Mammoth Mk II enroute.  Estimated ETA in 2 minutes...L   EVA: GDI援军已经到达. 猛犸机甲在路上, 预计2分钟后到达...%   EVA: Ghostalker lost, mission failed.%   EVA: 失去幽灵行者, 任务失败   EVA: Mammoth Mk II has arrived.   EVA: 猛犸机甲已经到达!   EVA: Mcneil lost, mission failed.(   EVA: 麦克尼尔失败了, 任务失败^   EVA: Penetrate their base, destroy that cargo car and retrieve the crate holding the crystals.K   EVA: 穿过他们的基地, 摧毁那辆货车, 取回装水晶的板条箱`   EVA: The bridge has been repaired and the train is making it's way to the Nod base in the south.;   EVA: 桥已经修好了火车正在往南边的Nod基地开X   EVA: The cargo car of that train contains the crate of crystals that you are to recover.F   EVA: 那列火车的货运车厢里有一箱水晶, 需要你去回收8   EVA: The crystals have been retrieved, mission complete.%   EVA: 水晶已经找到, 任务完成!   EVA: Umagon lost, mission failed."   EVA: 失去乌玛贡, 任务失败l   EVA: We are currently tracking the Nod train carrying the target cargo.  Intel states that the bridge is outR   EVA: 我们目前正在追踪Nod火车运载的目标货物. 情报显示桥断了"   Eye of the storm has been entered.   已进入风暴中心    Firestorm perimeter deactivated.   外围火焰风暴已关闭   First launcher deployed.   第一个发射器已经部署/   GDI Forces Spotted! Falling back to alert base.'   发现GDI部队! 回基地拉响警报!H   GDI Soldier: Shit, We're outnumbered! Return to base now and alert them.B   GDI士兵: 见鬼, 我们寡不敌众! 马上去基地拉响警报   GDI bullet train arriving.   GDI高速列车已抵达   GDI bullet train departing.   GDI高速列车已离开   GDI dropship detected.   探测到GDI运输机$   GDI forces spotted. Blow the bridge!   发现GDI部队. 把桥炸掉!   GDI has detected you.   GDI发现你了?   GDI is going after our extraction APC It must not be destroyed!9   GDI在追我们的运兵车, 绝对不能让它被干掉!*   GDI: Hurry Jake! They're right behind you!+   GDI: 快点, 杰克! 他们就在你后面!+   GDI: Jake, it's a trap! Get to the airbase!1   GDI: 杰克, 这是个陷阱! 快去空军基地!6   GDI: Jake, it's good to see...Hey! What are you doing?4   GDI: 杰克, 很高兴看到...嘿! 你在干什么?A   GDI: Jake, the transport will take 30 minutes to arrive. Hold on!<   GDI: 杰克, 运输机需要30分钟才能到达. 坚持住!6   GDI: Now watch the effectiveness against ground units.,   GDI: 现在看看对付地面单位的效果4   GDI: Patrol to base! Nod troops in area! Abort tour!@   GDI: 巡逻队返回基地! 发现Nod部队! 取消巡逻任务!5   GDI: The MM2 is equally deadly to air-based assaults.,   GDI: 猛犸机甲对空中攻击同样致命3   GDI: The MM2 is quite effective against structures.&   GDI: 猛犸机甲对建筑相当有效6   GDI: This concludes the Mammoth Mark II demonstration.&   GDI: 猛犸机甲的演示到此结束G   GDI: We've lost the beacon. Extraction time will be delayed 15 minutes.9   GDI: 我们失去了信标. 撤离时间将延迟15分钟M   Ghost Stalker: If you can get me onto that train, we can do some real damage!V   幽灵行者: 如果你能让我登上火车, 我们就能造成一些实质的伤害!"   Harvest the Tiberium to the north.   采集北方的泰伯利亚   Hassan Soldier: Hold them here!$   哈桑士兵: 把他们挡在这里!)   Hey! Where'd all those shiners come from?!   嘿! 这些闪光是从哪来的?:   Hey... over here! Help... Destroy these trucks to free us.@   嘿...这里! 帮帮我们...摧毁这些卡车, 放我们出来+   Holy $#!+ its Nod! I have to warn the base.%   见鬼! 是Nod! 我得去基地报告   ICBM destroyed!   已摧毁洲际弹道导弹!   ICBM launch detected.!   探测到洲际弹道导弹发射+   ICBMs destroyed! Philidephia out of danger.>   洲际弹道导弹被摧毁了! 费城空间站脱离了危险U   If your Tiberium Refinery is full, build Tiberium Silos to store the excess Tiberium.P   如果你的泰矿精炼厂满了, 建造泰矿储存仓来储存多余的泰矿   Kodiak destroyed!   科迪亚克被摧毁!   Kodiak in critical condition!   科迪亚克情况危急!   Kodiak under attack!   科迪亚克遭到攻击!   Laser Turrets! RUN FOR IT!   激光炮塔! 离它远点!   Launcher destroyed.   已摧毁发射器.9   Looks like they're going to ship it out via bullet train.$   看来他们要用火车运出去了5   Maximum efficiency for equipment can now be achieved.   设备已达到最大效率   Mission failed.   任务失败了!   Move quickly, before they see us.)   在他们看到我们之前, 赶紧行动   Mutant vermin detected.   发现变种害虫P   Mutants: Damn, their base has been cloaked. We must wait for them to uncloak it.H   变种人: 该死, 他们的基地隐形了, 我们得等他们漏出来5   Mutants: Hold a moment, while their fighters pass by.%   变种人: 等一下, 有敌人经过@   Mutants: Liars! GDI is trying to help us! You will die for this!F   变种人: 骗子! GDI是为了帮助我们! 你会为此付出代价!   Mutants: Okay, Go now.   变种人: 好了, 走吧N   Mutants: The charges are placed. We can get the laser wall down in 30 minutes.B   变种人: 炸药已安放. 我们能在30分钟内拆掉激光墙d   Mutants: The production facility has been located. Send in the reinforcements and let's finish this.N   变种人: 生产设备已经找到了. 派援军来, 让我们结束这一切4   Mutants: The wall is down - you are clear to attack!8   变种人: 激光墙已拆除, 你可以发动攻击了!D   New Objective: Get Ghost Stalker onto the train. Ghost must not die!=   新目标: 让幽灵行者登上火车. 记住, 他不能死!A   New secondary objective: Destroy primary AND secondary Nod bases.2   新次要目标: 摧毁Nod的主基地和次基地8   Nod ICBMs detected. To stop them, DESTROY the launchers.D   探测到Nod洲际弹道导弹. 摧毁导弹发射器以阻止他们f   Nod base is heavily guarded by lasers. Suggestion: destroying power plants to west may cause overload.a   Nod基地受到激光炮塔的严密保护. 建议: 摧毁西面的发电厂可使其电力超载X   Nod:  We can use these old units to our advantage.  Rerouting their control to you in 3,\   Nod: 我们可以利用这些老东西. 正在将它们的控制权转给你，3秒后完成I   Nod: All sensor arrays are down. Full area map generation dowloading now.C   Nod: 所有传感器阵列已瘫痪. 正在下载完整区域地图W   Nod: Commander, you have been provided with a direct satellite uplink for this mission.I   Nod: 指挥官, 本次任务已为你配备了直接的卫星上行链路]   Nod: Look to your radar now and you will see the three locations of the mobile sensor arrays.O   Nod: 现在看看你的雷达, 你会看到三个移动传感器阵列的位置8   Nod: Umagon has been detected in the northeast quadrant.    Nod: 在东北方发现乌玛贡1   Nod: Umagon has escaped. Your mission has failed.-   Nod: 乌玛贡已逃脱.你的任务失败了Z   Nod: Umagon has reached the GDI base and is moving to board the train leaving this region.F   Nod: 乌玛贡已到达GDI基地, 准备登上离开该地区的火车b   Nod: Umagon is moving to board the northern train which leaves the region. Her escape is imminent.=   Nod: 乌玛贡正准备登上北方的火车, 她要逃走了[   Nod: Umagon's dropship transport has arrived and she is moving to board the southern train.F   Nod: 乌玛贡的运输机已抵达, 她正准备登上南方的火车P   Nod: Umagon's dropship transport has been located and will arrive in 10 minutes.1   Nod: 乌玛贡的运输机将在10分钟后抵达9   Nod: Umagon's dropship transport will arrive in 1 minute.0   Nod: 乌玛贡的运输机将在1分钟后抵达:   Nod: Umagon's dropship transport will arrive in 5 minutes.0   Nod: 乌玛贡的运输机将在5分钟后抵达P   Note that your power is getting low. To get more power, build more Power Plants.c   请注意, 你的可用电力正在下降. 为了获得更多的电力, 请建造更多的发电厂[   Now get an engineer over here to fix this bridge and I will alert Hassan to their presence.M   现在找个工程师过来修理这座桥, 我将通知哈桑他们的位置   O.K.! You're clear to enter.   好的! 你可以进去了   Objective 1 complete.   目标一完成Z   Objective 1: Build a Tiberium Refinery and begin harvesting the Tiberium to the southeast.I   目标一: 建造一座泰矿精炼厂, 并开始在东南方开采泰矿7   Objective 1: Capture Hassan's T.V. station to the east.)   目标一: 占领东部哈桑的电视台8   Objective 1: Capture the GDI base before McNeil arrives.5   目标一: 在麦克尼尔到达之前占领GDI基地f   Objective 1: Capture the remaining GDI structures within this base to build a force to capture Tratos.^   目标一: 占领这个基地内剩余的GDI建筑, 并建立一支部队来抓捕特拉托斯I   Objective 1: Contact the mutants - try searching near the local hospital.G   目标一: 与变种人取得联系 - 尝试在当地医院附近搜索8   Objective 1: Deploy the ICBM launchers near the beacons.;   目标一: 在信标附近部署洲际弹道导弹发射器)   Objective 1: Destroy Nod missile complex.    目标一: 摧毁Nod导弹阵列(   Objective 1: Destroy all Nod structures.    目标一: 摧毁所有Nod建筑7   Objective 1: Destroy all chemical missile launch sites.,   目标一: 摧毁所有化学导弹发射台1   Objective 1: Destroy all of Hassan's elite guard.,   目标一: 摧毁哈桑所有的精锐卫队,   Objective 1: Destroy all the chemical tanks.&   目标一: 摧毁所有的化学储罐%   Objective 1: Destroy the supply base.   目标一: 摧毁补给基地B   Objective 1: Establish a base and build a Tiberium Waste Facility.&   目标一: 建造泰矿物质回收厂   Objective 1: Establish a base.   目标一: 建立基地$   Objective 1: Find and rescue Oxanna.)   目标一: 找到并营救奥克斯安娜>   Objective 1: Infiltrate the GDI Communication Upgrade Centers.    目标一: 渗透GDI通讯中心)   Objective 1: Locate and free the mutants.#   目标一: 定位并释放突变体.   Objective 1: Locate and secure the crash site.&   目标一: 定位并保护坠机现场8   Objective 1: Locate the abandoned Nod base to the north.)   目标一: 找到北部废弃的Nod基地N   Objective 1: Locate the crashed UFO and retrieve Kane's artifacts from inside.R   目标一: 找到坠毁的不明飞行物, 并从内部取回凯恩想要的东西*   Objective 1: Locate the old Temple of Nod.    目标一: 找到Nod的旧神殿%   Objective 1: Locate the toxin trucks.   目标一: 找到毒素卡车2   Objective 1: Plant C4 on all ten Nod power plants.(   目标一: 在所有Nod发电厂安装C4-   Objective 1: Protect the Kodiak at all costs./   目标一: 不惜一切代价保护科迪亚克3   Objective 1: Remove all Nod presence from the area.,   目标一: 清除该区域内所有Nod部队N   Objective 1: Spy on GDI comm center to learn the location of the weapons test.:   目标一: 潜入GDI通讯中心, 获取武器试验地点5   Objective 1: Stop the launch of the Tiberium Missile.)   目标一: 阻止泰伯利亚导弹发射   Objective 2 complete.   目标二完成6   Objective 2: Build a Barracks to create more infantry.,   目标二: 建造兵营来制造更多步兵%   Objective 2: Build the Temple of Nod.   目标二: 建造Nod神殿+   Objective 2: Capture Nod Technology Center.    目标二: 占领Nod技术中心$   Objective 2: Capture Vega's Pyramid.#   目标二: 占领维加的金字塔:   Objective 2: Capture the train station. DO NOT DESTROY IT!,   目标二: 占领火车站, 不要毁了它!7   Objective 2: Clear both ends of the tunnel to the west.&   目标二: 清除西边隧道的两头.   Objective 2: Commandeer a transport to escape.)   目标二: 抢占一辆运输车以逃离/   Objective 2: Destroy Hassan's elite guard base.,   目标二: 摧毁哈桑的精英卫队基地$   Objective 2: Destroy all Nod forces.    目标二: 摧毁所有Nod部队,   Objective 2: Destroy all five Nod SAM sites.,   目标二: 摧毁所有防空导弹发射台"   Objective 2: Destroy the GDI base.   目标二: 摧毁GDI基地;   Objective 2: Destroy the ICBMs targeted at the Philidephia.;   目标二: 摧毁针对费城空间站的洲际弹道导弹3   Objective 2: Destroy the Mammoth Mark II prototype.#   目标二: 摧毁猛犸机甲原型"   Objective 2: Destroy the Nod base.   目标二: 摧毁Nod基地I   Objective 2: Escort the toxin trucks past the GDI checkpoint to the east.8   目标二: 护送毒素卡车通过东部的GDI检查站(   Objective 2: Evacuate the Chameleon Spy.    目标二: 撤离变色龙间谍"   Objective 2: Evacuate the mutants.   目标二: 撤离变种人�   Objective 2: Now find the Mutant Headquarters and knock on their door (attack it!). This should convince Tratos to be sympathetic to our cause.u   目标二: 找到变种人总部并敲敲他们的门(攻击它!).这应该能说服特拉托斯加入我们的事业(   Objective 2: Remove the GDI trespassers.   目的二: 清除GDI入侵者/   Objective 2: Retrieve the cargo from the train.#   目标二: 从火车上取回货物@   Objective 2: To get production online build a Tiberium Refinery.1   目标二: 建设泰矿精炼厂, 使生产上线@   Objective 2: Use Toxin Soldiers to "convince" McNeil to join us.=   目标二: 利用毒素步兵"说服"麦克尼尔加入我们0   Objective 3: Destroy all Nod forces in the area.,   目标三: 摧毁该地区的所有Nod部队$   Objective 3: Destroy all Nod forces.    目标三: 摧毁所有Nod部队=   Objective 3: Get McNeil into the APC at the extraction point.5   目标三: 让麦克尼尔进入撤离点的运兵车7   Objective 3: Locate the research facility to the north.&   目标三: 找到北方的研究设施+   Objective 4: Destroy the research facility.   目标四: 摧毁研究设施'   Objective Reached: Civilians evacuated.   目标达成: 撤离平民!   Objective Reached: Mutants freed.   目标达成: 释放变种人   Objective Reached: Site secure   目标达成: 清除发射台.   Objective Reached: Technology Center captured.    目标达成: 占领技术中心7   Objective: Rescue captives from the prison to the east.&   目标: 营救东部监狱中的俘虏   One launcher remaining.   还剩一个发射器F   Orca Transport: Negative on extraction until SAM sites are eliminated!J   奥卡运输机: 在地对空导弹阵地未被清除前无法执行撤离9   Our cover is blown! Capture McNeil by any means possible!<   我们的身份暴露了! 尽一切可能抓住麦克尼尔!+   Oxanna is being moved to the main GDI base.3   奥克斯安娜正在被转移到GDI的主要基地   Oxanna located.   已找到奥克斯安娜   PEACE THROUGH POWER!   以力量实现和平!%   Perimeter secure. Deactivating alarm.   周边安全.关闭警报   Philidelphia in range.   空间站已在射程内2   Power levels are low. Construct more Power Plants./   电力水平低. 需要建造更多的发电厂   Power overload in progress...   电力过载...:   Prevent the train from departing and retreive the Tacitus.&   阻止火车出发, 并取回塔西佗1   Proceed to the next Communication Upgrade Center.!   前往下一个通信升级中心*   Proceed with Tiberium Missile destruction.*   继续执行泰伯利亚导弹摧毁任务   Pull over for inspection!   靠边接受检查!)   Reentering ion storm, caution is advised.3   重新进入离子风暴区域，建议小心行事   SCROOGE!
   小气鬼!   STOP THAT TRAIN!   停下那列火车!   Second launcher deployed.   第二个发射器已部署<   She is boarding a train bound for the GDI base in the south.-   她正在登上开往南部GDI基地的火车M   Sir! I believe there is an old GDI base near. It could be worth looking into.F   长官! 我发现附近有一个废弃的GDI基地, 可能值得调查8   Sir! The Tacitus is gone. Vega's men must've grabbed it.:   长官! 塔西佗不见了, 肯定被维加的人抢走了p   Solomon: Change of plans - We have verified Vega's presence in the pyramid. CAPTURE the pyramid with Vega alive.m   所罗门: 计划有变 - 我们已经证实了维加在金字塔中的存在. 逮捕维加并占领金字塔*   Sound the Alarm! Slavik's Forces are here!*   拉响警报! 斯拉维克的军队来了!   Special objective complete.   特殊目标完成0   Stand and Identify yourself in the name of Kane.,   以凯恩之名, 停下并表明你的身份    Stand forward and be recognized!   站过来, 接受身份识别!1   Stop! Don't Shoot! I was forced to work for them.4   停下! 不要开枪! 我是被迫为他们工作的-   Storm abating. Commence attack on Nod forces.#   风暴减弱, 开始攻击Nod部队   Supplies found.   已找到补给   Tacitus has been acquired.   已被获取塔西佗@   Take out this sentry post and I will show you their nearby base.;   摧毁这个哨兵岗, 我会带你去他们附近的基地   Thanks for the help!   谢谢你的帮助!;   Thanks! We can use the supplies.  I'll go gather my people.:   谢谢! 我们正需要这些补给, 我去叫我的人来$   The Philadelphia has been destroyed!   费城空间站被摧毁了!%   The Philidelphia has left ICBM range.3   费城空间站已脱离洲际弹道导弹的射程.   The Philidelphia is passing within ICBM Range.3   费城空间站正进入洲际弹道导弹射程内   The Temple is under attack!   神殿遭到攻击!@   The temple has been discovered, NOW DESTROY the GDI trespassers.2   神殿已被发现, 现在摧毁所有GDI入侵者,   The traitors are coming, destroy the bridge!   叛徒来了, 摧毁这座桥!0   They are sending a transmission to Sarajevo now.'   他们正在向萨拉热窝发送信号,   Third launcher deployed. Objective complete./   第三个发射装置已经部署. 目标完成   This map is under redesign.!   这张地图正在重新设计中   Tiberium Missile launched.   泰伯利亚导弹已发射   Tiberium lifeform detected.   检测到泰伯生命体"   Tiberium waste convoy approaching.!   泰矿物质运输车正在靠近A   To build or train left-click on the icons located in the sidebar.8   要建造或生产, 请左键点击侧边栏中的图标V   To deploy a vehicle select it, place the cursor over the vehicle and left-click on it.Q   要部署载具, 先选择它, 然后将光标移至载具上, 最后左键点击N   To repair a bridge, send an engineer into the repair hut near the bridge base.J   要修复桥梁, 请派遣一名工程师进入桥基附近的修理工棚c   To repair a structure left-click on the wrench icon in the sidebar and left-click on the structure.X   要修复建筑, 先左键点击侧边栏的扳手图标, 然后左键点击目标建筑   Transport has arrived.   运输机已抵达   Transport lost.   失去运输机;   Tratos: Fight them my children, for the fate of our people.E   特拉托斯: 族人们, 为了我们种族的命运, 与他们战斗V   Tratos: You have killed enough of my children, take me and be done with this violence.N   特拉托斯: 你们已经杀了我太多族人, 带我走吧, 结束这暴力   Two launchers remaining.   还剩两个发射器   UFO crash sight located.   发现不明飞行物信号   Umagon: My people are nearby.    乌玛贡: 我的人就在附近5   Umagon: My people are waiting somewhere to the north.,   乌玛贡: 我的族人在北方某处等着6   Use the Weedeater units to harvest the Tiberium veins.-   使用除草机单位采集泰伯利亚矿脉1   Warning: Mission critical structure under attack.&   警告: 关键任务建造受到攻击,   Warning: Mission critical unit under attack.&   警告: 关键任务单位受到攻击X   We have Hassan pinned and ready to be brought in Commander Slavick. Orders are complete.7   我们已将哈桑围困, 正在抓捕, 任务已完成*   We have to get this to Tratos immediately.-   我们必须马上把这个交给特拉托斯7   We should rendezvous with the rescue team to the south.'   我们应该和南方的救援队会合   We will help.   我们会提供帮助^   We've been touched by the spirit hand of Kane, and are ready to serve the technology of peace.G   我们已接受凯恩神灵之手的感召, 准备为和平科技效力?   What's the E.T.A. on that M.C.V.? This UFO gives me the creeps.>   那台基地车还有多久到? 这个飞船让我毛骨悚然d   You have been provided with 2 Artillery units. Good hunting, reinforcements will be arriving soon...C   你已得到两台炮兵单位. 狩猎愉快, 增援很快到达...=   Your venture has been quite unsuccessful, to state the least.)   不委婉地说, 你的行动相当失败7   and we may hit the train before they repair the bridge.3   如果我们能在他们修好桥之前拦下火车C   to the South. Penetrate the bases defenses and retrieve that cargo.,   到南方. 穿透基地防御并取回货物ui    $  '   (Use -1 to signify an unlimited supply)   (使用-1表示无限补给)   1 on 1   1 v 1   2 on 2   2 v 2   < Back   < 返回	   AI Level:	   AI级别:
   AI Players   电脑玩家   AI Players:   电脑玩家:   Abort   放弃   Abort Mission   放弃任务   Accept   接受   Accessability:   可访问性:   Action Message   动作资讯   Add   添加   Allies Allowed   已允许结盟   Allies allowed   已允许结盟   Allow incoming pages       Allow others to find me   允许别人查找我   Answer   应答   Assign   分配   Available Servers   可用服务器   Ban a user from your channel$   禁止一个用户进入你的频道   Bases   基地
   BattleClan
   BattleClan   BattleClan Tournament   BattleClan 锦标赛   BattleClan Tournament Webpage   BattleClan 锦标赛网页   Baud:
   波特率:   Better   更好	   Birthdate   生日   Bridges Destroyable   可摧毁桥梁   Button 3   按钮 3   Call Waiting:   等待呼叫:
   Cameo Text   图标文本   Cancel   取消	   Category:   类别:   Channel Password:   频道密码:   Cities:   城市:Z   Click OK to keep this display mode or wait and your old display settings will be restored.P   单击"确定"以保持此显示模式, 或者等待恢复您的旧显示设置.   Cliffs:   悬崖:   Color:   颜色:	   Commands:   命令:
   Connection   连接   Continue   继续   Crates	   板条箱   Create Random Map   建立随机地图   Create a new chat channel:   创建新的聊天频道:   Credits	   制作组   Credits:   资金:   Current shortcut:   当前快捷键:   Currently assigned to:   当前分配到:   Custom	   自定义   Customize Keyboard   自定义键盘   DELETE   删除   Data Compression   数据压缩   Debug   调试   Default   默认   Delete   删除   Delete Game   删除游戏
   Delete Map   删除地图   Description   描述   Description:   描述:   Destination Network:   目标网络:   Details:   细节:   Dial   拨号
   Difficulty   难度
   Disconnect   断开连接   Disconnects   断开连接   Display   显示   Display Options:   显示选项:!   Do you want to abort the mission?   你想放弃当前任务吗?   Down   下   Downloading patch   正在下载补丁   Dropship Loadout Limits   运输船装卸限制   Dropship Unit Limit   运输船单位限制   Edit   编辑4   Email address:           (Please double check this!)'   电子邮件地址:     (双击这个!)   Environment:   环境:   Error Correction   误差修正   Exit   退出	   Exit Game   退出游戏   Faster   更快   Filter bad language   过滤不良语言   Find   查找   Find a game   查找游戏   Find/Page another user   查找/分页其他用户	   Firestorm   火焰风暴
   Fog Of War   战争迷雾   Game Controls   游戏控制   Game Settings   游戏设置
   Game Speed   游戏速度   Game Speed:   游戏速度:	   Game Type   游戏类型   Games   游戏   Games:   游戏:   Get a Westwood Online login   获取Westwood在线登录   Go to the BattleClan webpage   转到BattleClan网页   Go!   开始!   Harder   更难   Harvester Truce   采矿车休战   Help   帮助   Higher   更高   Hills:   山丘:   Host Location   主机位置?   I would like to receive the Westwood Online newsletter by Email;   我想通过电子邮件接收Westwood网络的时事通讯	   IPX (Lan)   IPX(局域网)   IPX Options
   IPX 选项   Ignore a user   忽略一个用户   Init String   初始化字符串   Internet	   互联网   Internet Game Controls   网络游戏控制   Intro / Sneak Peek   简介/先睹为快
   Ion Storms   离子风暴   Join   加入   Join Battle Clan   加入BattleClan   Keyboard   键盘   Kick a user from your channel!   把一个用户踢出你的频道
   Kill Limit   击杀限制   LOAD   加载   Ladder Rank of Host   房主排名   Ladder:   阶梯:	   Lifeforms	   生命体   Load   加载	   Load Game   加载游戏   Load Map   加载地图   Load Mission   加载任务	   Location:   地区:   Losses   损失	   Main Menu	   主菜单   Map   地图   Map Height:   地图高度:
   Map Width:   地图宽度:   Map:   地图:   Max   最大   Max Ping to Host   到主机的最大Ping   Max Players   最大玩家数   Min   最小   Mission   任务   Modem / Serial   调制解调器 / 串口   Multi Engineer   多位工程师   Multiplay Map   多人地图   Multiplayer Game   多人游戏   Multiplayer Map   多人游戏地图   Music Volume:   音乐音量:   Name   名称   Name:   名称:   Network   网络   Network Card:   网卡:   New   新建   New Account	   新帐号   New Campaign	   新战役   Next >   继续 >	   Nickname:   昵称:   No   否   None   无
   Null Modem   调制解调器   Number:   数量:   OK   确定   Official   官方	   Opponent:   对手:   Options   选项   Options Menu   选项菜单   Page   页	   Page Clan       Parent's Email address:   家长的电子邮件地址:	   Password:   密码:   Person to find or page:   要查找或分页的人:
   Phone List   电话列表   Phone Number:   电话号码   Phonebook Entry   电话簿条目   Play   播放
   Play music   播放音乐   Player   玩家   Player 1   玩家 1   Player 2   玩家 2   Player 3   玩家 3   Player 4   玩家 4   Player 5   玩家 5   Player 6   玩家 6   Player 7   玩家 7   Player 8   玩家 8   Player Tournament Webpage   玩家锦标赛网页   Players   玩家   Players:   玩家:3   Please visit our website at http://www.westwood.com3   请访问我我们的网页 http://www.westwood.com   Points   点   Port:   端口:   Press new shortcut key:   按下新的快捷键:   Preview   预览   Preview Map   预览地图	   Progress1   进度1
   Pulse Dial   脉冲拨号   Quit   退出   Random   随机   Rank   排名   Re-Deployable MCV   可重新部署MCV   Re-enter Password:   重新输入密码:   Refresh Channel List   刷新频道列表   Refresh Channels   刷新频道   Repeat   重复	   Reset All   全部重置   Resolution Modes   分辨率模式   Restart   重新开始   Restate Briefing   重述简报   Resume Mission   恢复任务   SAVE   保存   Save   保存	   Save Game   保存游戏   Save Map   保存地图   Scroll Coasting   惯性滚动   Scroll Rate   滚动速率   Scroll Rate:   滚动速率:   Search:   搜索:   Select Campaign:   选择战役:   Select Game Type   选择游戏类型   Select Multiplayer Game   选择多人游戏   Select Multiplayer Map   选择多人游戏地图   Selected Game Details   选定游戏详情   Serial Settings   串口设置   Server:
   服务器:   Set Location   设置位置   Settings   设置	   Settings:   设置:
   Short Game   快速游戏   Show All   全部显示   Show all games in my lobby!   在我的大厅展示所有游戏   Shuffle   随机   Side:   阵营:   Sidebar Text   侧边栏文本   Skirmish	   遭遇战   Slider1   滑块1   Slider2   滑块2   Slider3   滑块3   Slider4   滑块4   Slider5   滑块5   Slider6   滑块6   Socket Number:   Socket 号码:   Sound   声音   Sound Options   声音选项   Sound Volume:   音量:   Squad   分组   Standard   标准   Stop   停止   Store login   登录店铺    Stretch movies to fit resolution   拉伸电影以适应分辨率   Surprise Me   随机生成   Target Lines	   目标线
   Tech Level   科技等级   Tech Level:   科技等级:   Text to send:   要发送的文本:   Tiberian Sun   泰伯利亚之日   Tiberian Sun (Original)   泰伯利亚之日 (原版)'   Tiberian Sun Has Encountered Difficulty!   泰伯利亚之日遇到了问题K   Tiberian Sun has encountered a problem.
See the file DEBUG.TXT for details.N   泰伯利亚之日遇到了一个问题.
详细信息请参见DEBUG.TXT文件..   Tiberian Sun has encountered an internal error-   泰伯利亚之日遇到了一个内部错误   Tiberium Amount:   泰矿数量:   Tiberium Fields:
   泰矿田:
   Time Limit   时间限制   Time Remaining:   剩余时间:
   Time Stamp   时间   Time of Day:   时间:	   Tone Dial   按键式拨号   Tooltips   工具提示
   Tournament	   锦标赛   Transitions   过渡   UDP (Internet)   UDP (互联网)
   Unit Count   单位数量   Unit Count:   单位数量:	   Unit Name   单位名称   Unknown	   未知的   Up   上   Users:   用户:   Vegetation:   植被:
   Veinholes:
   脉络孔:   View the privacy policy   查看隐私政策   View the tournament ladder   查看锦标赛天梯   Visual Details   视觉细节   Visual Details:   视觉细节:   Voice Volume:   语音音量:   Waiting for a response   等待响应   Water:   水体:   Westwood Online options   Westwood在线选项   Wins   获胜�   World Domination Tour games use your Battle Clan affiliation to determine which side you are fighting for.  If you do not wish to join a Battle Clan, select which side you wish to fight for.�   世界统治之旅使用你的Battle Clan隶属关系来确定你为哪一方而战. 如果你不想加入Battle Clan, 请选择你的阵营.   World Domination! (Internet)   统治世界! (互联网)   Yes   是�   Yes, EA/Westwood can share the information I have provided with other companies so they can notify me of new products and special offers.j   是的, EA/Westwood可以与其他公司分享我提供的信息, 以便他们通知我新产品和促销.   Your Color:   你的颜色:   Your Location   你的位置
   Your Name:   你的名字:
   Your Side:   你的阵营:%   Your password must be 8 letters long.&   您的密码长度必须为8个字母.#   and is unable to continue normally.   并且无法正常继续.-   for the latest updates and technical support.%   获取最新的更新和技术支持.